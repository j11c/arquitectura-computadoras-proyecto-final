-------------------------------------------------------------------------------
--
-- Company : Universidad Miguel Hernandez
-- Engineer: joshi
-- 
-- Create Date:    30/11/2025 10:21:36
-- Project Name:   computadora_didactica
-- Module Name:    computadora_didactica_tb.vhd
-- Description:
--
-- Additional Comments:
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;  -- Para std_logic
use IEEE.numeric_std.all;     -- Para signed, unsigned

entity computadora_didactica_tb is
end    computadora_didactica_tb;

architecture Testbench of computadora_didactica_tb is

   -- Component Declaration for the Unit Under Test (UUT)
   component computadora_didactica
	port( 
		clk		: in std_logic;
		entrada : in std_logic_vector(11 downto 0);
		salida	: out std_logic_vector(11 downto 0);
		halted	: out std_logic
	);
   end component;

   -- Select an architecture if needed (default is last one analyzed).
   --for uut: computadora_didactica use entity WORK.computadora_didactica(arq1);

   -- Inputs/Outputs
   signal entrada, salida : std_logic_vector(11 downto 0) := x"000";
   signal halted : std_logic := '0';

   -- Clock (uncomment if needed)
   -- Sustituir <clock> por el nombre de puerto apropiado
   signal   clk : std_logic := '0';
   constant clock_period : time := 50 ns;
   signal   clock_on : boolean := true;

begin

   -- Instantiate the Unit Under Test (UUT)
   uut: computadora_didactica port map ( 
		clk => clk,
		entrada => entrada,
		salida => salida,
		halted => halted
   );

-- Clock process (uncomment if needed)
-- Descomentar en caso de requerir senial de reloj
-- Sustituir <clock> por el nombre de puerto apropiado
clock_process : process
begin
   while (clock_on) loop
      clk <= '0';
      wait for clock_period/2;
      clk <= '1';
      wait for clock_period/2;
   end loop;
   --assert (false) report ("Finished") severity error;
   -- Wait forever
   wait;
 end process;

-- Stimulus process
stim_proc: process
begin
   -- hold reset state for 100 ns
   wait for 100 ns;

   ---------------------------------------------------------
   -- insert stimulus here
   ---------------------------------------------------------

   -- Test case 1
   -- ... Asignaciones a seniales de entrada ...
   wait for 1000 ns;
   -- assert (<condition>) report "Error case 1" severity error;

   -- Test case 2
   -- ... Asignaciones a seniales de entrada ...
   wait for 100 ns;
   -- assert (<condition>) report "Error case 2" severity error;

   -- Stop clock
   clock_on <= false;
   -- Wait forever
   wait;

end process;

end Testbench;
