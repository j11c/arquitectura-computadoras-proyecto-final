-------------------------------------------------------------------------------
--
-- Company : Universidad Miguel Hernandez
-- Engineer: joshi
-- 
-- Create Date:    20/11/2025 09:37:07
-- Project Name:   memoriaPrograma
-- Module Name:    memoriaPrograma.vhd
-- Description:
--
-- Additional Comments:
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;  -- Para std_logic
use IEEE.numeric_std.all;     -- Para unsigned

entity memoriaPrograma is
	port( 
		addr : in  std_logic_vector(9 downto 0);
        data : out std_logic_vector(9 downto 0)
	);
end memoriaPrograma;

architecture arq1 of memoriaPrograma is
	
	type mem_type is array (0 to 1023) of std_logic_vector(9 downto 0);

	constant ROM : mem_type := (
"1001110100", -- linea 1 / direccion 0x000 (0)
"0000000001", -- linea 2 / direccion 0x001 (1)
"1001110000", -- linea 3 / direccion 0x002 (2)
"0000000010", -- linea 4 / direccion 0x003 (3)
"1000000001", -- linea 5 / direccion 0x004 (4)
"1101110000", -- linea 6 / direccion 0x005 (5)
"0000001001", -- linea 7 / direccion 0x006 (6)
"0001110000", -- linea 8 / direccion 0x007 (7)
"0000001010", -- linea 9 / direccion 0x008 (8)
"1100100000", -- linea 10 / direccion 0x009 (9)
"1111000000", -- linea 11 / direccion 0x00A (10)
"0000000000", -- linea 12 / direccion 0x00B (11) (NOP)
"0000000000", -- linea 13 / direccion 0x00C (12) (NOP)
"0000000000", -- linea 14 / direccion 0x00D (13) (NOP)
"0000000000", -- linea 15 / direccion 0x00E (14) (NOP)
"0000000000", -- linea 16 / direccion 0x00F (15) (NOP)
    "0000000000", -- linea 17 / direccion 0x010 (16) (NOP)
    "0000000000", -- linea 18 / direccion 0x011 (17) (NOP)
    "0000000000", -- linea 19 / direccion 0x012 (18) (NOP)
    "0000000000", -- linea 20 / direccion 0x013 (19) (NOP)
    "0000000000", -- linea 21 / direccion 0x014 (20) (NOP)
    "0000000000", -- linea 22 / direccion 0x015 (21) (NOP)
    "0000000000", -- linea 23 / direccion 0x016 (22) (NOP)
    "0000000000", -- linea 24 / direccion 0x017 (23) (NOP)
    "0000000000", -- linea 25 / direccion 0x018 (24) (NOP)
    "0000000000", -- linea 26 / direccion 0x019 (25) (NOP)
    "0000000000", -- linea 27 / direccion 0x01A (26) (NOP)
    "0000000000", -- linea 28 / direccion 0x01B (27) (NOP)
    "0000000000", -- linea 29 / direccion 0x01C (28) (NOP)
    "0000000000", -- linea 30 / direccion 0x01D (29) (NOP)
    "0000000000", -- linea 31 / direccion 0x01E (30) (NOP)
    "0000000000", -- linea 32 / direccion 0x01F (31) (NOP)
    "0000000000", -- linea 33 / direccion 0x020 (32) (NOP)
    "0000000000", -- linea 34 / direccion 0x021 (33) (NOP)
    "0000000000", -- linea 35 / direccion 0x022 (34) (NOP)
    "0000000000", -- linea 36 / direccion 0x023 (35) (NOP)
    "0000000000", -- linea 37 / direccion 0x024 (36) (NOP)
    "0000000000", -- linea 38 / direccion 0x025 (37) (NOP)
    "0000000000", -- linea 39 / direccion 0x026 (38) (NOP)
    "0000000000", -- linea 40 / direccion 0x027 (39) (NOP)
    "0000000000", -- linea 41 / direccion 0x028 (40) (NOP)
    "0000000000", -- linea 42 / direccion 0x029 (41) (NOP)
    "0000000000", -- linea 43 / direccion 0x02A (42) (NOP)
    "0000000000", -- linea 44 / direccion 0x02B (43) (NOP)
    "0000000000", -- linea 45 / direccion 0x02C (44) (NOP)
    "0000000000", -- linea 46 / direccion 0x02D (45) (NOP)
    "0000000000", -- linea 47 / direccion 0x02E (46) (NOP)
    "0000000000", -- linea 48 / direccion 0x02F (47) (NOP)
    "0000000000", -- linea 49 / direccion 0x030 (48) (NOP)
    "0000000000", -- linea 50 / direccion 0x031 (49) (NOP)
    "0000000000", -- linea 51 / direccion 0x032 (50) (NOP)
    "0000000000", -- linea 52 / direccion 0x033 (51) (NOP)
    "0000000000", -- linea 53 / direccion 0x034 (52) (NOP)
    "0000000000", -- linea 54 / direccion 0x035 (53) (NOP)
    "0000000000", -- linea 55 / direccion 0x036 (54) (NOP)
    "0000000000", -- linea 56 / direccion 0x037 (55) (NOP)
    "0000000000", -- linea 57 / direccion 0x038 (56) (NOP)
    "0000000000", -- linea 58 / direccion 0x039 (57) (NOP)
    "0000000000", -- linea 59 / direccion 0x03A (58) (NOP)
    "0000000000", -- linea 60 / direccion 0x03B (59) (NOP)
    "0000000000", -- linea 61 / direccion 0x03C (60) (NOP)
    "0000000000", -- linea 62 / direccion 0x03D (61) (NOP)
    "0000000000", -- linea 63 / direccion 0x03E (62) (NOP)
    "0000000000", -- linea 64 / direccion 0x03F (63) (NOP)
    "0000000000", -- linea 65 / direccion 0x040 (64) (NOP)
    "0000000000", -- linea 66 / direccion 0x041 (65) (NOP)
    "0000000000", -- linea 67 / direccion 0x042 (66) (NOP)
    "0000000000", -- linea 68 / direccion 0x043 (67) (NOP)
    "0000000000", -- linea 69 / direccion 0x044 (68) (NOP)
    "0000000000", -- linea 70 / direccion 0x045 (69) (NOP)
    "0000000000", -- linea 71 / direccion 0x046 (70) (NOP)
    "0000000000", -- linea 72 / direccion 0x047 (71) (NOP)
    "0000000000", -- linea 73 / direccion 0x048 (72) (NOP)
    "0000000000", -- linea 74 / direccion 0x049 (73) (NOP)
    "0000000000", -- linea 75 / direccion 0x04A (74) (NOP)
    "0000000000", -- linea 76 / direccion 0x04B (75) (NOP)
    "0000000000", -- linea 77 / direccion 0x04C (76) (NOP)
    "0000000000", -- linea 78 / direccion 0x04D (77) (NOP)
    "0000000000", -- linea 79 / direccion 0x04E (78) (NOP)
    "0000000000", -- linea 80 / direccion 0x04F (79) (NOP)
    "0000000000", -- linea 81 / direccion 0x050 (80) (NOP)
    "0000000000", -- linea 82 / direccion 0x051 (81) (NOP)
    "0000000000", -- linea 83 / direccion 0x052 (82) (NOP)
    "0000000000", -- linea 84 / direccion 0x053 (83) (NOP)
    "0000000000", -- linea 85 / direccion 0x054 (84) (NOP)
    "0000000000", -- linea 86 / direccion 0x055 (85) (NOP)
    "0000000000", -- linea 87 / direccion 0x056 (86) (NOP)
    "0000000000", -- linea 88 / direccion 0x057 (87) (NOP)
    "0000000000", -- linea 89 / direccion 0x058 (88) (NOP)
    "0000000000", -- linea 90 / direccion 0x059 (89) (NOP)
    "0000000000", -- linea 91 / direccion 0x05A (90) (NOP)
    "0000000000", -- linea 92 / direccion 0x05B (91) (NOP)
    "0000000000", -- linea 93 / direccion 0x05C (92) (NOP)
    "0000000000", -- linea 94 / direccion 0x05D (93) (NOP)
    "0000000000", -- linea 95 / direccion 0x05E (94) (NOP)
    "0000000000", -- linea 96 / direccion 0x05F (95) (NOP)
    "0000000000", -- linea 97 / direccion 0x060 (96) (NOP)
    "0000000000", -- linea 98 / direccion 0x061 (97) (NOP)
    "0000000000", -- linea 99 / direccion 0x062 (98) (NOP)
    "0000000000", -- linea 100 / direccion 0x063 (99) (NOP)
    "0000000000", -- linea 101 / direccion 0x064 (100) (NOP)
    "0000000000", -- linea 102 / direccion 0x065 (101) (NOP)
    "0000000000", -- linea 103 / direccion 0x066 (102) (NOP)
    "0000000000", -- linea 104 / direccion 0x067 (103) (NOP)
    "0000000000", -- linea 105 / direccion 0x068 (104) (NOP)
    "0000000000", -- linea 106 / direccion 0x069 (105) (NOP)
    "0000000000", -- linea 107 / direccion 0x06A (106) (NOP)
    "0000000000", -- linea 108 / direccion 0x06B (107) (NOP)
    "0000000000", -- linea 109 / direccion 0x06C (108) (NOP)
    "0000000000", -- linea 110 / direccion 0x06D (109) (NOP)
    "0000000000", -- linea 111 / direccion 0x06E (110) (NOP)
    "0000000000", -- linea 112 / direccion 0x06F (111) (NOP)
    "0000000000", -- linea 113 / direccion 0x070 (112) (NOP)
    "0000000000", -- linea 114 / direccion 0x071 (113) (NOP)
    "0000000000", -- linea 115 / direccion 0x072 (114) (NOP)
    "0000000000", -- linea 116 / direccion 0x073 (115) (NOP)
    "0000000000", -- linea 117 / direccion 0x074 (116) (NOP)
    "0000000000", -- linea 118 / direccion 0x075 (117) (NOP)
    "0000000000", -- linea 119 / direccion 0x076 (118) (NOP)
    "0000000000", -- linea 120 / direccion 0x077 (119) (NOP)
    "0000000000", -- linea 121 / direccion 0x078 (120) (NOP)
    "0000000000", -- linea 122 / direccion 0x079 (121) (NOP)
    "0000000000", -- linea 123 / direccion 0x07A (122) (NOP)
    "0000000000", -- linea 124 / direccion 0x07B (123) (NOP)
    "0000000000", -- linea 125 / direccion 0x07C (124) (NOP)
    "0000000000", -- linea 126 / direccion 0x07D (125) (NOP)
    "0000000000", -- linea 127 / direccion 0x07E (126) (NOP)
    "0000000000", -- linea 128 / direccion 0x07F (127) (NOP)
    "0000000000", -- linea 129 / direccion 0x080 (128) (NOP)
    "0000000000", -- linea 130 / direccion 0x081 (129) (NOP)
    "0000000000", -- linea 131 / direccion 0x082 (130) (NOP)
    "0000000000", -- linea 132 / direccion 0x083 (131) (NOP)
    "0000000000", -- linea 133 / direccion 0x084 (132) (NOP)
    "0000000000", -- linea 134 / direccion 0x085 (133) (NOP)
    "0000000000", -- linea 135 / direccion 0x086 (134) (NOP)
    "0000000000", -- linea 136 / direccion 0x087 (135) (NOP)
    "0000000000", -- linea 137 / direccion 0x088 (136) (NOP)
    "0000000000", -- linea 138 / direccion 0x089 (137) (NOP)
    "0000000000", -- linea 139 / direccion 0x08A (138) (NOP)
    "0000000000", -- linea 140 / direccion 0x08B (139) (NOP)
    "0000000000", -- linea 141 / direccion 0x08C (140) (NOP)
    "0000000000", -- linea 142 / direccion 0x08D (141) (NOP)
    "0000000000", -- linea 143 / direccion 0x08E (142) (NOP)
    "0000000000", -- linea 144 / direccion 0x08F (143) (NOP)
    "0000000000", -- linea 145 / direccion 0x090 (144) (NOP)
    "0000000000", -- linea 146 / direccion 0x091 (145) (NOP)
    "0000000000", -- linea 147 / direccion 0x092 (146) (NOP)
    "0000000000", -- linea 148 / direccion 0x093 (147) (NOP)
    "0000000000", -- linea 149 / direccion 0x094 (148) (NOP)
    "0000000000", -- linea 150 / direccion 0x095 (149) (NOP)
    "0000000000", -- linea 151 / direccion 0x096 (150) (NOP)
    "0000000000", -- linea 152 / direccion 0x097 (151) (NOP)
    "0000000000", -- linea 153 / direccion 0x098 (152) (NOP)
    "0000000000", -- linea 154 / direccion 0x099 (153) (NOP)
    "0000000000", -- linea 155 / direccion 0x09A (154) (NOP)
    "0000000000", -- linea 156 / direccion 0x09B (155) (NOP)
    "0000000000", -- linea 157 / direccion 0x09C (156) (NOP)
    "0000000000", -- linea 158 / direccion 0x09D (157) (NOP)
    "0000000000", -- linea 159 / direccion 0x09E (158) (NOP)
    "0000000000", -- linea 160 / direccion 0x09F (159) (NOP)
    "0000000000", -- linea 161 / direccion 0x0A0 (160) (NOP)
    "0000000000", -- linea 162 / direccion 0x0A1 (161) (NOP)
    "0000000000", -- linea 163 / direccion 0x0A2 (162) (NOP)
    "0000000000", -- linea 164 / direccion 0x0A3 (163) (NOP)
    "0000000000", -- linea 165 / direccion 0x0A4 (164) (NOP)
    "0000000000", -- linea 166 / direccion 0x0A5 (165) (NOP)
    "0000000000", -- linea 167 / direccion 0x0A6 (166) (NOP)
    "0000000000", -- linea 168 / direccion 0x0A7 (167) (NOP)
    "0000000000", -- linea 169 / direccion 0x0A8 (168) (NOP)
    "0000000000", -- linea 170 / direccion 0x0A9 (169) (NOP)
    "0000000000", -- linea 171 / direccion 0x0AA (170) (NOP)
    "0000000000", -- linea 172 / direccion 0x0AB (171) (NOP)
    "0000000000", -- linea 173 / direccion 0x0AC (172) (NOP)
    "0000000000", -- linea 174 / direccion 0x0AD (173) (NOP)
    "0000000000", -- linea 175 / direccion 0x0AE (174) (NOP)
    "0000000000", -- linea 176 / direccion 0x0AF (175) (NOP)
    "0000000000", -- linea 177 / direccion 0x0B0 (176) (NOP)
    "0000000000", -- linea 178 / direccion 0x0B1 (177) (NOP)
    "0000000000", -- linea 179 / direccion 0x0B2 (178) (NOP)
    "0000000000", -- linea 180 / direccion 0x0B3 (179) (NOP)
    "0000000000", -- linea 181 / direccion 0x0B4 (180) (NOP)
    "0000000000", -- linea 182 / direccion 0x0B5 (181) (NOP)
    "0000000000", -- linea 183 / direccion 0x0B6 (182) (NOP)
    "0000000000", -- linea 184 / direccion 0x0B7 (183) (NOP)
    "0000000000", -- linea 185 / direccion 0x0B8 (184) (NOP)
    "0000000000", -- linea 186 / direccion 0x0B9 (185) (NOP)
    "0000000000", -- linea 187 / direccion 0x0BA (186) (NOP)
    "0000000000", -- linea 188 / direccion 0x0BB (187) (NOP)
    "0000000000", -- linea 189 / direccion 0x0BC (188) (NOP)
    "0000000000", -- linea 190 / direccion 0x0BD (189) (NOP)
    "0000000000", -- linea 191 / direccion 0x0BE (190) (NOP)
    "0000000000", -- linea 192 / direccion 0x0BF (191) (NOP)
    "0000000000", -- linea 193 / direccion 0x0C0 (192) (NOP)
    "0000000000", -- linea 194 / direccion 0x0C1 (193) (NOP)
    "0000000000", -- linea 195 / direccion 0x0C2 (194) (NOP)
    "0000000000", -- linea 196 / direccion 0x0C3 (195) (NOP)
    "0000000000", -- linea 197 / direccion 0x0C4 (196) (NOP)
    "0000000000", -- linea 198 / direccion 0x0C5 (197) (NOP)
    "0000000000", -- linea 199 / direccion 0x0C6 (198) (NOP)
    "0000000000", -- linea 200 / direccion 0x0C7 (199) (NOP)
    "0000000000", -- linea 201 / direccion 0x0C8 (200) (NOP)
    "0000000000", -- linea 202 / direccion 0x0C9 (201) (NOP)
    "0000000000", -- linea 203 / direccion 0x0CA (202) (NOP)
    "0000000000", -- linea 204 / direccion 0x0CB (203) (NOP)
    "0000000000", -- linea 205 / direccion 0x0CC (204) (NOP)
    "0000000000", -- linea 206 / direccion 0x0CD (205) (NOP)
    "0000000000", -- linea 207 / direccion 0x0CE (206) (NOP)
    "0000000000", -- linea 208 / direccion 0x0CF (207) (NOP)
    "0000000000", -- linea 209 / direccion 0x0D0 (208) (NOP)
    "0000000000", -- linea 210 / direccion 0x0D1 (209) (NOP)
    "0000000000", -- linea 211 / direccion 0x0D2 (210) (NOP)
    "0000000000", -- linea 212 / direccion 0x0D3 (211) (NOP)
    "0000000000", -- linea 213 / direccion 0x0D4 (212) (NOP)
    "0000000000", -- linea 214 / direccion 0x0D5 (213) (NOP)
    "0000000000", -- linea 215 / direccion 0x0D6 (214) (NOP)
    "0000000000", -- linea 216 / direccion 0x0D7 (215) (NOP)
    "0000000000", -- linea 217 / direccion 0x0D8 (216) (NOP)
    "0000000000", -- linea 218 / direccion 0x0D9 (217) (NOP)
    "0000000000", -- linea 219 / direccion 0x0DA (218) (NOP)
    "0000000000", -- linea 220 / direccion 0x0DB (219) (NOP)
    "0000000000", -- linea 221 / direccion 0x0DC (220) (NOP)
    "0000000000", -- linea 222 / direccion 0x0DD (221) (NOP)
    "0000000000", -- linea 223 / direccion 0x0DE (222) (NOP)
    "0000000000", -- linea 224 / direccion 0x0DF (223) (NOP)
    "0000000000", -- linea 225 / direccion 0x0E0 (224) (NOP)
    "0000000000", -- linea 226 / direccion 0x0E1 (225) (NOP)
    "0000000000", -- linea 227 / direccion 0x0E2 (226) (NOP)
    "0000000000", -- linea 228 / direccion 0x0E3 (227) (NOP)
    "0000000000", -- linea 229 / direccion 0x0E4 (228) (NOP)
    "0000000000", -- linea 230 / direccion 0x0E5 (229) (NOP)
    "0000000000", -- linea 231 / direccion 0x0E6 (230) (NOP)
    "0000000000", -- linea 232 / direccion 0x0E7 (231) (NOP)
    "0000000000", -- linea 233 / direccion 0x0E8 (232) (NOP)
    "0000000000", -- linea 234 / direccion 0x0E9 (233) (NOP)
    "0000000000", -- linea 235 / direccion 0x0EA (234) (NOP)
    "0000000000", -- linea 236 / direccion 0x0EB (235) (NOP)
    "0000000000", -- linea 237 / direccion 0x0EC (236) (NOP)
    "0000000000", -- linea 238 / direccion 0x0ED (237) (NOP)
    "0000000000", -- linea 239 / direccion 0x0EE (238) (NOP)
    "0000000000", -- linea 240 / direccion 0x0EF (239) (NOP)
    "0000000000", -- linea 241 / direccion 0x0F0 (240) (NOP)
    "0000000000", -- linea 242 / direccion 0x0F1 (241) (NOP)
    "0000000000", -- linea 243 / direccion 0x0F2 (242) (NOP)
    "0000000000", -- linea 244 / direccion 0x0F3 (243) (NOP)
    "0000000000", -- linea 245 / direccion 0x0F4 (244) (NOP)
    "0000000000", -- linea 246 / direccion 0x0F5 (245) (NOP)
    "0000000000", -- linea 247 / direccion 0x0F6 (246) (NOP)
    "0000000000", -- linea 248 / direccion 0x0F7 (247) (NOP)
    "0000000000", -- linea 249 / direccion 0x0F8 (248) (NOP)
    "0000000000", -- linea 250 / direccion 0x0F9 (249) (NOP)
    "0000000000", -- linea 251 / direccion 0x0FA (250) (NOP)
    "0000000000", -- linea 252 / direccion 0x0FB (251) (NOP)
    "0000000000", -- linea 253 / direccion 0x0FC (252) (NOP)
    "0000000000", -- linea 254 / direccion 0x0FD (253) (NOP)
    "0000000000", -- linea 255 / direccion 0x0FE (254) (NOP)
    "0000000000", -- linea 256 / direccion 0x0FF (255) (NOP)
    "0000000000", -- linea 257 / direccion 0x100 (256) (NOP)
    "0000000000", -- linea 258 / direccion 0x101 (257) (NOP)
    "0000000000", -- linea 259 / direccion 0x102 (258) (NOP)
    "0000000000", -- linea 260 / direccion 0x103 (259) (NOP)
    "0000000000", -- linea 261 / direccion 0x104 (260) (NOP)
    "0000000000", -- linea 262 / direccion 0x105 (261) (NOP)
    "0000000000", -- linea 263 / direccion 0x106 (262) (NOP)
    "0000000000", -- linea 264 / direccion 0x107 (263) (NOP)
    "0000000000", -- linea 265 / direccion 0x108 (264) (NOP)
    "0000000000", -- linea 266 / direccion 0x109 (265) (NOP)
    "0000000000", -- linea 267 / direccion 0x10A (266) (NOP)
    "0000000000", -- linea 268 / direccion 0x10B (267) (NOP)
    "0000000000", -- linea 269 / direccion 0x10C (268) (NOP)
    "0000000000", -- linea 270 / direccion 0x10D (269) (NOP)
    "0000000000", -- linea 271 / direccion 0x10E (270) (NOP)
    "0000000000", -- linea 272 / direccion 0x10F (271) (NOP)
    "0000000000", -- linea 273 / direccion 0x110 (272) (NOP)
    "0000000000", -- linea 274 / direccion 0x111 (273) (NOP)
    "0000000000", -- linea 275 / direccion 0x112 (274) (NOP)
    "0000000000", -- linea 276 / direccion 0x113 (275) (NOP)
    "0000000000", -- linea 277 / direccion 0x114 (276) (NOP)
    "0000000000", -- linea 278 / direccion 0x115 (277) (NOP)
    "0000000000", -- linea 279 / direccion 0x116 (278) (NOP)
    "0000000000", -- linea 280 / direccion 0x117 (279) (NOP)
    "0000000000", -- linea 281 / direccion 0x118 (280) (NOP)
    "0000000000", -- linea 282 / direccion 0x119 (281) (NOP)
    "0000000000", -- linea 283 / direccion 0x11A (282) (NOP)
    "0000000000", -- linea 284 / direccion 0x11B (283) (NOP)
    "0000000000", -- linea 285 / direccion 0x11C (284) (NOP)
    "0000000000", -- linea 286 / direccion 0x11D (285) (NOP)
    "0000000000", -- linea 287 / direccion 0x11E (286) (NOP)
    "0000000000", -- linea 288 / direccion 0x11F (287) (NOP)
    "0000000000", -- linea 289 / direccion 0x120 (288) (NOP)
    "0000000000", -- linea 290 / direccion 0x121 (289) (NOP)
    "0000000000", -- linea 291 / direccion 0x122 (290) (NOP)
    "0000000000", -- linea 292 / direccion 0x123 (291) (NOP)
    "0000000000", -- linea 293 / direccion 0x124 (292) (NOP)
    "0000000000", -- linea 294 / direccion 0x125 (293) (NOP)
    "0000000000", -- linea 295 / direccion 0x126 (294) (NOP)
    "0000000000", -- linea 296 / direccion 0x127 (295) (NOP)
    "0000000000", -- linea 297 / direccion 0x128 (296) (NOP)
    "0000000000", -- linea 298 / direccion 0x129 (297) (NOP)
    "0000000000", -- linea 299 / direccion 0x12A (298) (NOP)
    "0000000000", -- linea 300 / direccion 0x12B (299) (NOP)
    "0000000000", -- linea 301 / direccion 0x12C (300) (NOP)
    "0000000000", -- linea 302 / direccion 0x12D (301) (NOP)
    "0000000000", -- linea 303 / direccion 0x12E (302) (NOP)
    "0000000000", -- linea 304 / direccion 0x12F (303) (NOP)
    "0000000000", -- linea 305 / direccion 0x130 (304) (NOP)
    "0000000000", -- linea 306 / direccion 0x131 (305) (NOP)
    "0000000000", -- linea 307 / direccion 0x132 (306) (NOP)
    "0000000000", -- linea 308 / direccion 0x133 (307) (NOP)
    "0000000000", -- linea 309 / direccion 0x134 (308) (NOP)
    "0000000000", -- linea 310 / direccion 0x135 (309) (NOP)
    "0000000000", -- linea 311 / direccion 0x136 (310) (NOP)
    "0000000000", -- linea 312 / direccion 0x137 (311) (NOP)
    "0000000000", -- linea 313 / direccion 0x138 (312) (NOP)
    "0000000000", -- linea 314 / direccion 0x139 (313) (NOP)
    "0000000000", -- linea 315 / direccion 0x13A (314) (NOP)
    "0000000000", -- linea 316 / direccion 0x13B (315) (NOP)
    "0000000000", -- linea 317 / direccion 0x13C (316) (NOP)
    "0000000000", -- linea 318 / direccion 0x13D (317) (NOP)
    "0000000000", -- linea 319 / direccion 0x13E (318) (NOP)
    "0000000000", -- linea 320 / direccion 0x13F (319) (NOP)
    "0000000000", -- linea 321 / direccion 0x140 (320) (NOP)
    "0000000000", -- linea 322 / direccion 0x141 (321) (NOP)
    "0000000000", -- linea 323 / direccion 0x142 (322) (NOP)
    "0000000000", -- linea 324 / direccion 0x143 (323) (NOP)
    "0000000000", -- linea 325 / direccion 0x144 (324) (NOP)
    "0000000000", -- linea 326 / direccion 0x145 (325) (NOP)
    "0000000000", -- linea 327 / direccion 0x146 (326) (NOP)
    "0000000000", -- linea 328 / direccion 0x147 (327) (NOP)
    "0000000000", -- linea 329 / direccion 0x148 (328) (NOP)
    "0000000000", -- linea 330 / direccion 0x149 (329) (NOP)
    "0000000000", -- linea 331 / direccion 0x14A (330) (NOP)
    "0000000000", -- linea 332 / direccion 0x14B (331) (NOP)
    "0000000000", -- linea 333 / direccion 0x14C (332) (NOP)
    "0000000000", -- linea 334 / direccion 0x14D (333) (NOP)
    "0000000000", -- linea 335 / direccion 0x14E (334) (NOP)
    "0000000000", -- linea 336 / direccion 0x14F (335) (NOP)
    "0000000000", -- linea 337 / direccion 0x150 (336) (NOP)
    "0000000000", -- linea 338 / direccion 0x151 (337) (NOP)
    "0000000000", -- linea 339 / direccion 0x152 (338) (NOP)
    "0000000000", -- linea 340 / direccion 0x153 (339) (NOP)
    "0000000000", -- linea 341 / direccion 0x154 (340) (NOP)
    "0000000000", -- linea 342 / direccion 0x155 (341) (NOP)
    "0000000000", -- linea 343 / direccion 0x156 (342) (NOP)
    "0000000000", -- linea 344 / direccion 0x157 (343) (NOP)
    "0000000000", -- linea 345 / direccion 0x158 (344) (NOP)
    "0000000000", -- linea 346 / direccion 0x159 (345) (NOP)
    "0000000000", -- linea 347 / direccion 0x15A (346) (NOP)
    "0000000000", -- linea 348 / direccion 0x15B (347) (NOP)
    "0000000000", -- linea 349 / direccion 0x15C (348) (NOP)
    "0000000000", -- linea 350 / direccion 0x15D (349) (NOP)
    "0000000000", -- linea 351 / direccion 0x15E (350) (NOP)
    "0000000000", -- linea 352 / direccion 0x15F (351) (NOP)
    "0000000000", -- linea 353 / direccion 0x160 (352) (NOP)
    "0000000000", -- linea 354 / direccion 0x161 (353) (NOP)
    "0000000000", -- linea 355 / direccion 0x162 (354) (NOP)
    "0000000000", -- linea 356 / direccion 0x163 (355) (NOP)
    "0000000000", -- linea 357 / direccion 0x164 (356) (NOP)
    "0000000000", -- linea 358 / direccion 0x165 (357) (NOP)
    "0000000000", -- linea 359 / direccion 0x166 (358) (NOP)
    "0000000000", -- linea 360 / direccion 0x167 (359) (NOP)
    "0000000000", -- linea 361 / direccion 0x168 (360) (NOP)
    "0000000000", -- linea 362 / direccion 0x169 (361) (NOP)
    "0000000000", -- linea 363 / direccion 0x16A (362) (NOP)
    "0000000000", -- linea 364 / direccion 0x16B (363) (NOP)
    "0000000000", -- linea 365 / direccion 0x16C (364) (NOP)
    "0000000000", -- linea 366 / direccion 0x16D (365) (NOP)
    "0000000000", -- linea 367 / direccion 0x16E (366) (NOP)
    "0000000000", -- linea 368 / direccion 0x16F (367) (NOP)
    "0000000000", -- linea 369 / direccion 0x170 (368) (NOP)
    "0000000000", -- linea 370 / direccion 0x171 (369) (NOP)
    "0000000000", -- linea 371 / direccion 0x172 (370) (NOP)
    "0000000000", -- linea 372 / direccion 0x173 (371) (NOP)
    "0000000000", -- linea 373 / direccion 0x174 (372) (NOP)
    "0000000000", -- linea 374 / direccion 0x175 (373) (NOP)
    "0000000000", -- linea 375 / direccion 0x176 (374) (NOP)
    "0000000000", -- linea 376 / direccion 0x177 (375) (NOP)
    "0000000000", -- linea 377 / direccion 0x178 (376) (NOP)
    "0000000000", -- linea 378 / direccion 0x179 (377) (NOP)
    "0000000000", -- linea 379 / direccion 0x17A (378) (NOP)
    "0000000000", -- linea 380 / direccion 0x17B (379) (NOP)
    "0000000000", -- linea 381 / direccion 0x17C (380) (NOP)
    "0000000000", -- linea 382 / direccion 0x17D (381) (NOP)
    "0000000000", -- linea 383 / direccion 0x17E (382) (NOP)
    "0000000000", -- linea 384 / direccion 0x17F (383) (NOP)
    "0000000000", -- linea 385 / direccion 0x180 (384) (NOP)
    "0000000000", -- linea 386 / direccion 0x181 (385) (NOP)
    "0000000000", -- linea 387 / direccion 0x182 (386) (NOP)
    "0000000000", -- linea 388 / direccion 0x183 (387) (NOP)
    "0000000000", -- linea 389 / direccion 0x184 (388) (NOP)
    "0000000000", -- linea 390 / direccion 0x185 (389) (NOP)
    "0000000000", -- linea 391 / direccion 0x186 (390) (NOP)
    "0000000000", -- linea 392 / direccion 0x187 (391) (NOP)
    "0000000000", -- linea 393 / direccion 0x188 (392) (NOP)
    "0000000000", -- linea 394 / direccion 0x189 (393) (NOP)
    "0000000000", -- linea 395 / direccion 0x18A (394) (NOP)
    "0000000000", -- linea 396 / direccion 0x18B (395) (NOP)
    "0000000000", -- linea 397 / direccion 0x18C (396) (NOP)
    "0000000000", -- linea 398 / direccion 0x18D (397) (NOP)
    "0000000000", -- linea 399 / direccion 0x18E (398) (NOP)
    "0000000000", -- linea 400 / direccion 0x18F (399) (NOP)
    "0000000000", -- linea 401 / direccion 0x190 (400) (NOP)
    "0000000000", -- linea 402 / direccion 0x191 (401) (NOP)
    "0000000000", -- linea 403 / direccion 0x192 (402) (NOP)
    "0000000000", -- linea 404 / direccion 0x193 (403) (NOP)
    "0000000000", -- linea 405 / direccion 0x194 (404) (NOP)
    "0000000000", -- linea 406 / direccion 0x195 (405) (NOP)
    "0000000000", -- linea 407 / direccion 0x196 (406) (NOP)
    "0000000000", -- linea 408 / direccion 0x197 (407) (NOP)
    "0000000000", -- linea 409 / direccion 0x198 (408) (NOP)
    "0000000000", -- linea 410 / direccion 0x199 (409) (NOP)
    "0000000000", -- linea 411 / direccion 0x19A (410) (NOP)
    "0000000000", -- linea 412 / direccion 0x19B (411) (NOP)
    "0000000000", -- linea 413 / direccion 0x19C (412) (NOP)
    "0000000000", -- linea 414 / direccion 0x19D (413) (NOP)
    "0000000000", -- linea 415 / direccion 0x19E (414) (NOP)
    "0000000000", -- linea 416 / direccion 0x19F (415) (NOP)
    "0000000000", -- linea 417 / direccion 0x1A0 (416) (NOP)
    "0000000000", -- linea 418 / direccion 0x1A1 (417) (NOP)
    "0000000000", -- linea 419 / direccion 0x1A2 (418) (NOP)
    "0000000000", -- linea 420 / direccion 0x1A3 (419) (NOP)
    "0000000000", -- linea 421 / direccion 0x1A4 (420) (NOP)
    "0000000000", -- linea 422 / direccion 0x1A5 (421) (NOP)
    "0000000000", -- linea 423 / direccion 0x1A6 (422) (NOP)
    "0000000000", -- linea 424 / direccion 0x1A7 (423) (NOP)
    "0000000000", -- linea 425 / direccion 0x1A8 (424) (NOP)
    "0000000000", -- linea 426 / direccion 0x1A9 (425) (NOP)
    "0000000000", -- linea 427 / direccion 0x1AA (426) (NOP)
    "0000000000", -- linea 428 / direccion 0x1AB (427) (NOP)
    "0000000000", -- linea 429 / direccion 0x1AC (428) (NOP)
    "0000000000", -- linea 430 / direccion 0x1AD (429) (NOP)
    "0000000000", -- linea 431 / direccion 0x1AE (430) (NOP)
    "0000000000", -- linea 432 / direccion 0x1AF (431) (NOP)
    "0000000000", -- linea 433 / direccion 0x1B0 (432) (NOP)
    "0000000000", -- linea 434 / direccion 0x1B1 (433) (NOP)
    "0000000000", -- linea 435 / direccion 0x1B2 (434) (NOP)
    "0000000000", -- linea 436 / direccion 0x1B3 (435) (NOP)
    "0000000000", -- linea 437 / direccion 0x1B4 (436) (NOP)
    "0000000000", -- linea 438 / direccion 0x1B5 (437) (NOP)
    "0000000000", -- linea 439 / direccion 0x1B6 (438) (NOP)
    "0000000000", -- linea 440 / direccion 0x1B7 (439) (NOP)
    "0000000000", -- linea 441 / direccion 0x1B8 (440) (NOP)
    "0000000000", -- linea 442 / direccion 0x1B9 (441) (NOP)
    "0000000000", -- linea 443 / direccion 0x1BA (442) (NOP)
    "0000000000", -- linea 444 / direccion 0x1BB (443) (NOP)
    "0000000000", -- linea 445 / direccion 0x1BC (444) (NOP)
    "0000000000", -- linea 446 / direccion 0x1BD (445) (NOP)
    "0000000000", -- linea 447 / direccion 0x1BE (446) (NOP)
    "0000000000", -- linea 448 / direccion 0x1BF (447) (NOP)
    "0000000000", -- linea 449 / direccion 0x1C0 (448) (NOP)
    "0000000000", -- linea 450 / direccion 0x1C1 (449) (NOP)
    "0000000000", -- linea 451 / direccion 0x1C2 (450) (NOP)
    "0000000000", -- linea 452 / direccion 0x1C3 (451) (NOP)
    "0000000000", -- linea 453 / direccion 0x1C4 (452) (NOP)
    "0000000000", -- linea 454 / direccion 0x1C5 (453) (NOP)
    "0000000000", -- linea 455 / direccion 0x1C6 (454) (NOP)
    "0000000000", -- linea 456 / direccion 0x1C7 (455) (NOP)
    "0000000000", -- linea 457 / direccion 0x1C8 (456) (NOP)
    "0000000000", -- linea 458 / direccion 0x1C9 (457) (NOP)
    "0000000000", -- linea 459 / direccion 0x1CA (458) (NOP)
    "0000000000", -- linea 460 / direccion 0x1CB (459) (NOP)
    "0000000000", -- linea 461 / direccion 0x1CC (460) (NOP)
    "0000000000", -- linea 462 / direccion 0x1CD (461) (NOP)
    "0000000000", -- linea 463 / direccion 0x1CE (462) (NOP)
    "0000000000", -- linea 464 / direccion 0x1CF (463) (NOP)
    "0000000000", -- linea 465 / direccion 0x1D0 (464) (NOP)
    "0000000000", -- linea 466 / direccion 0x1D1 (465) (NOP)
    "0000000000", -- linea 467 / direccion 0x1D2 (466) (NOP)
    "0000000000", -- linea 468 / direccion 0x1D3 (467) (NOP)
    "0000000000", -- linea 469 / direccion 0x1D4 (468) (NOP)
    "0000000000", -- linea 470 / direccion 0x1D5 (469) (NOP)
    "0000000000", -- linea 471 / direccion 0x1D6 (470) (NOP)
    "0000000000", -- linea 472 / direccion 0x1D7 (471) (NOP)
    "0000000000", -- linea 473 / direccion 0x1D8 (472) (NOP)
    "0000000000", -- linea 474 / direccion 0x1D9 (473) (NOP)
    "0000000000", -- linea 475 / direccion 0x1DA (474) (NOP)
    "0000000000", -- linea 476 / direccion 0x1DB (475) (NOP)
    "0000000000", -- linea 477 / direccion 0x1DC (476) (NOP)
    "0000000000", -- linea 478 / direccion 0x1DD (477) (NOP)
    "0000000000", -- linea 479 / direccion 0x1DE (478) (NOP)
    "0000000000", -- linea 480 / direccion 0x1DF (479) (NOP)
    "0000000000", -- linea 481 / direccion 0x1E0 (480) (NOP)
    "0000000000", -- linea 482 / direccion 0x1E1 (481) (NOP)
    "0000000000", -- linea 483 / direccion 0x1E2 (482) (NOP)
    "0000000000", -- linea 484 / direccion 0x1E3 (483) (NOP)
    "0000000000", -- linea 485 / direccion 0x1E4 (484) (NOP)
    "0000000000", -- linea 486 / direccion 0x1E5 (485) (NOP)
    "0000000000", -- linea 487 / direccion 0x1E6 (486) (NOP)
    "0000000000", -- linea 488 / direccion 0x1E7 (487) (NOP)
    "0000000000", -- linea 489 / direccion 0x1E8 (488) (NOP)
    "0000000000", -- linea 490 / direccion 0x1E9 (489) (NOP)
    "0000000000", -- linea 491 / direccion 0x1EA (490) (NOP)
    "0000000000", -- linea 492 / direccion 0x1EB (491) (NOP)
    "0000000000", -- linea 493 / direccion 0x1EC (492) (NOP)
    "0000000000", -- linea 494 / direccion 0x1ED (493) (NOP)
    "0000000000", -- linea 495 / direccion 0x1EE (494) (NOP)
    "0000000000", -- linea 496 / direccion 0x1EF (495) (NOP)
    "0000000000", -- linea 497 / direccion 0x1F0 (496) (NOP)
    "0000000000", -- linea 498 / direccion 0x1F1 (497) (NOP)
    "0000000000", -- linea 499 / direccion 0x1F2 (498) (NOP)
    "0000000000", -- linea 500 / direccion 0x1F3 (499) (NOP)
    "0000000000", -- linea 501 / direccion 0x1F4 (500) (NOP)
    "0000000000", -- linea 502 / direccion 0x1F5 (501) (NOP)
    "0000000000", -- linea 503 / direccion 0x1F6 (502) (NOP)
    "0000000000", -- linea 504 / direccion 0x1F7 (503) (NOP)
    "0000000000", -- linea 505 / direccion 0x1F8 (504) (NOP)
    "0000000000", -- linea 506 / direccion 0x1F9 (505) (NOP)
    "0000000000", -- linea 507 / direccion 0x1FA (506) (NOP)
    "0000000000", -- linea 508 / direccion 0x1FB (507) (NOP)
    "0000000000", -- linea 509 / direccion 0x1FC (508) (NOP)
    "0000000000", -- linea 510 / direccion 0x1FD (509) (NOP)
    "0000000000", -- linea 511 / direccion 0x1FE (510) (NOP)
    "0000000000", -- linea 512 / direccion 0x1FF (511) (NOP)
    "0000000000", -- linea 513 / direccion 0x200 (512) (NOP)
    "0000000000", -- linea 514 / direccion 0x201 (513) (NOP)
    "0000000000", -- linea 515 / direccion 0x202 (514) (NOP)
    "0000000000", -- linea 516 / direccion 0x203 (515) (NOP)
    "0000000000", -- linea 517 / direccion 0x204 (516) (NOP)
    "0000000000", -- linea 518 / direccion 0x205 (517) (NOP)
    "0000000000", -- linea 519 / direccion 0x206 (518) (NOP)
    "0000000000", -- linea 520 / direccion 0x207 (519) (NOP)
    "0000000000", -- linea 521 / direccion 0x208 (520) (NOP)
    "0000000000", -- linea 522 / direccion 0x209 (521) (NOP)
    "0000000000", -- linea 523 / direccion 0x20A (522) (NOP)
    "0000000000", -- linea 524 / direccion 0x20B (523) (NOP)
    "0000000000", -- linea 525 / direccion 0x20C (524) (NOP)
    "0000000000", -- linea 526 / direccion 0x20D (525) (NOP)
    "0000000000", -- linea 527 / direccion 0x20E (526) (NOP)
    "0000000000", -- linea 528 / direccion 0x20F (527) (NOP)
    "0000000000", -- linea 529 / direccion 0x210 (528) (NOP)
    "0000000000", -- linea 530 / direccion 0x211 (529) (NOP)
    "0000000000", -- linea 531 / direccion 0x212 (530) (NOP)
    "0000000000", -- linea 532 / direccion 0x213 (531) (NOP)
    "0000000000", -- linea 533 / direccion 0x214 (532) (NOP)
    "0000000000", -- linea 534 / direccion 0x215 (533) (NOP)
    "0000000000", -- linea 535 / direccion 0x216 (534) (NOP)
    "0000000000", -- linea 536 / direccion 0x217 (535) (NOP)
    "0000000000", -- linea 537 / direccion 0x218 (536) (NOP)
    "0000000000", -- linea 538 / direccion 0x219 (537) (NOP)
    "0000000000", -- linea 539 / direccion 0x21A (538) (NOP)
    "0000000000", -- linea 540 / direccion 0x21B (539) (NOP)
    "0000000000", -- linea 541 / direccion 0x21C (540) (NOP)
    "0000000000", -- linea 542 / direccion 0x21D (541) (NOP)
    "0000000000", -- linea 543 / direccion 0x21E (542) (NOP)
    "0000000000", -- linea 544 / direccion 0x21F (543) (NOP)
    "0000000000", -- linea 545 / direccion 0x220 (544) (NOP)
    "0000000000", -- linea 546 / direccion 0x221 (545) (NOP)
    "0000000000", -- linea 547 / direccion 0x222 (546) (NOP)
    "0000000000", -- linea 548 / direccion 0x223 (547) (NOP)
    "0000000000", -- linea 549 / direccion 0x224 (548) (NOP)
    "0000000000", -- linea 550 / direccion 0x225 (549) (NOP)
    "0000000000", -- linea 551 / direccion 0x226 (550) (NOP)
    "0000000000", -- linea 552 / direccion 0x227 (551) (NOP)
    "0000000000", -- linea 553 / direccion 0x228 (552) (NOP)
    "0000000000", -- linea 554 / direccion 0x229 (553) (NOP)
    "0000000000", -- linea 555 / direccion 0x22A (554) (NOP)
    "0000000000", -- linea 556 / direccion 0x22B (555) (NOP)
    "0000000000", -- linea 557 / direccion 0x22C (556) (NOP)
    "0000000000", -- linea 558 / direccion 0x22D (557) (NOP)
    "0000000000", -- linea 559 / direccion 0x22E (558) (NOP)
    "0000000000", -- linea 560 / direccion 0x22F (559) (NOP)
    "0000000000", -- linea 561 / direccion 0x230 (560) (NOP)
    "0000000000", -- linea 562 / direccion 0x231 (561) (NOP)
    "0000000000", -- linea 563 / direccion 0x232 (562) (NOP)
    "0000000000", -- linea 564 / direccion 0x233 (563) (NOP)
    "0000000000", -- linea 565 / direccion 0x234 (564) (NOP)
    "0000000000", -- linea 566 / direccion 0x235 (565) (NOP)
    "0000000000", -- linea 567 / direccion 0x236 (566) (NOP)
    "0000000000", -- linea 568 / direccion 0x237 (567) (NOP)
    "0000000000", -- linea 569 / direccion 0x238 (568) (NOP)
    "0000000000", -- linea 570 / direccion 0x239 (569) (NOP)
    "0000000000", -- linea 571 / direccion 0x23A (570) (NOP)
    "0000000000", -- linea 572 / direccion 0x23B (571) (NOP)
    "0000000000", -- linea 573 / direccion 0x23C (572) (NOP)
    "0000000000", -- linea 574 / direccion 0x23D (573) (NOP)
    "0000000000", -- linea 575 / direccion 0x23E (574) (NOP)
    "0000000000", -- linea 576 / direccion 0x23F (575) (NOP)
    "0000000000", -- linea 577 / direccion 0x240 (576) (NOP)
    "0000000000", -- linea 578 / direccion 0x241 (577) (NOP)
    "0000000000", -- linea 579 / direccion 0x242 (578) (NOP)
    "0000000000", -- linea 580 / direccion 0x243 (579) (NOP)
    "0000000000", -- linea 581 / direccion 0x244 (580) (NOP)
    "0000000000", -- linea 582 / direccion 0x245 (581) (NOP)
    "0000000000", -- linea 583 / direccion 0x246 (582) (NOP)
    "0000000000", -- linea 584 / direccion 0x247 (583) (NOP)
    "0000000000", -- linea 585 / direccion 0x248 (584) (NOP)
    "0000000000", -- linea 586 / direccion 0x249 (585) (NOP)
    "0000000000", -- linea 587 / direccion 0x24A (586) (NOP)
    "0000000000", -- linea 588 / direccion 0x24B (587) (NOP)
    "0000000000", -- linea 589 / direccion 0x24C (588) (NOP)
    "0000000000", -- linea 590 / direccion 0x24D (589) (NOP)
    "0000000000", -- linea 591 / direccion 0x24E (590) (NOP)
    "0000000000", -- linea 592 / direccion 0x24F (591) (NOP)
    "0000000000", -- linea 593 / direccion 0x250 (592) (NOP)
    "0000000000", -- linea 594 / direccion 0x251 (593) (NOP)
    "0000000000", -- linea 595 / direccion 0x252 (594) (NOP)
    "0000000000", -- linea 596 / direccion 0x253 (595) (NOP)
    "0000000000", -- linea 597 / direccion 0x254 (596) (NOP)
    "0000000000", -- linea 598 / direccion 0x255 (597) (NOP)
    "0000000000", -- linea 599 / direccion 0x256 (598) (NOP)
    "0000000000", -- linea 600 / direccion 0x257 (599) (NOP)
    "0000000000", -- linea 601 / direccion 0x258 (600) (NOP)
    "0000000000", -- linea 602 / direccion 0x259 (601) (NOP)
    "0000000000", -- linea 603 / direccion 0x25A (602) (NOP)
    "0000000000", -- linea 604 / direccion 0x25B (603) (NOP)
    "0000000000", -- linea 605 / direccion 0x25C (604) (NOP)
    "0000000000", -- linea 606 / direccion 0x25D (605) (NOP)
    "0000000000", -- linea 607 / direccion 0x25E (606) (NOP)
    "0000000000", -- linea 608 / direccion 0x25F (607) (NOP)
    "0000000000", -- linea 609 / direccion 0x260 (608) (NOP)
    "0000000000", -- linea 610 / direccion 0x261 (609) (NOP)
    "0000000000", -- linea 611 / direccion 0x262 (610) (NOP)
    "0000000000", -- linea 612 / direccion 0x263 (611) (NOP)
    "0000000000", -- linea 613 / direccion 0x264 (612) (NOP)
    "0000000000", -- linea 614 / direccion 0x265 (613) (NOP)
    "0000000000", -- linea 615 / direccion 0x266 (614) (NOP)
    "0000000000", -- linea 616 / direccion 0x267 (615) (NOP)
    "0000000000", -- linea 617 / direccion 0x268 (616) (NOP)
    "0000000000", -- linea 618 / direccion 0x269 (617) (NOP)
    "0000000000", -- linea 619 / direccion 0x26A (618) (NOP)
    "0000000000", -- linea 620 / direccion 0x26B (619) (NOP)
    "0000000000", -- linea 621 / direccion 0x26C (620) (NOP)
    "0000000000", -- linea 622 / direccion 0x26D (621) (NOP)
    "0000000000", -- linea 623 / direccion 0x26E (622) (NOP)
    "0000000000", -- linea 624 / direccion 0x26F (623) (NOP)
    "0000000000", -- linea 625 / direccion 0x270 (624) (NOP)
    "0000000000", -- linea 626 / direccion 0x271 (625) (NOP)
    "0000000000", -- linea 627 / direccion 0x272 (626) (NOP)
    "0000000000", -- linea 628 / direccion 0x273 (627) (NOP)
    "0000000000", -- linea 629 / direccion 0x274 (628) (NOP)
    "0000000000", -- linea 630 / direccion 0x275 (629) (NOP)
    "0000000000", -- linea 631 / direccion 0x276 (630) (NOP)
    "0000000000", -- linea 632 / direccion 0x277 (631) (NOP)
    "0000000000", -- linea 633 / direccion 0x278 (632) (NOP)
    "0000000000", -- linea 634 / direccion 0x279 (633) (NOP)
    "0000000000", -- linea 635 / direccion 0x27A (634) (NOP)
    "0000000000", -- linea 636 / direccion 0x27B (635) (NOP)
    "0000000000", -- linea 637 / direccion 0x27C (636) (NOP)
    "0000000000", -- linea 638 / direccion 0x27D (637) (NOP)
    "0000000000", -- linea 639 / direccion 0x27E (638) (NOP)
    "0000000000", -- linea 640 / direccion 0x27F (639) (NOP)
    "0000000000", -- linea 641 / direccion 0x280 (640) (NOP)
    "0000000000", -- linea 642 / direccion 0x281 (641) (NOP)
    "0000000000", -- linea 643 / direccion 0x282 (642) (NOP)
    "0000000000", -- linea 644 / direccion 0x283 (643) (NOP)
    "0000000000", -- linea 645 / direccion 0x284 (644) (NOP)
    "0000000000", -- linea 646 / direccion 0x285 (645) (NOP)
    "0000000000", -- linea 647 / direccion 0x286 (646) (NOP)
    "0000000000", -- linea 648 / direccion 0x287 (647) (NOP)
    "0000000000", -- linea 649 / direccion 0x288 (648) (NOP)
    "0000000000", -- linea 650 / direccion 0x289 (649) (NOP)
    "0000000000", -- linea 651 / direccion 0x28A (650) (NOP)
    "0000000000", -- linea 652 / direccion 0x28B (651) (NOP)
    "0000000000", -- linea 653 / direccion 0x28C (652) (NOP)
    "0000000000", -- linea 654 / direccion 0x28D (653) (NOP)
    "0000000000", -- linea 655 / direccion 0x28E (654) (NOP)
    "0000000000", -- linea 656 / direccion 0x28F (655) (NOP)
    "0000000000", -- linea 657 / direccion 0x290 (656) (NOP)
    "0000000000", -- linea 658 / direccion 0x291 (657) (NOP)
    "0000000000", -- linea 659 / direccion 0x292 (658) (NOP)
    "0000000000", -- linea 660 / direccion 0x293 (659) (NOP)
    "0000000000", -- linea 661 / direccion 0x294 (660) (NOP)
    "0000000000", -- linea 662 / direccion 0x295 (661) (NOP)
    "0000000000", -- linea 663 / direccion 0x296 (662) (NOP)
    "0000000000", -- linea 664 / direccion 0x297 (663) (NOP)
    "0000000000", -- linea 665 / direccion 0x298 (664) (NOP)
    "0000000000", -- linea 666 / direccion 0x299 (665) (NOP)
    "0000000000", -- linea 667 / direccion 0x29A (666) (NOP)
    "0000000000", -- linea 668 / direccion 0x29B (667) (NOP)
    "0000000000", -- linea 669 / direccion 0x29C (668) (NOP)
    "0000000000", -- linea 670 / direccion 0x29D (669) (NOP)
    "0000000000", -- linea 671 / direccion 0x29E (670) (NOP)
    "0000000000", -- linea 672 / direccion 0x29F (671) (NOP)
    "0000000000", -- linea 673 / direccion 0x2A0 (672) (NOP)
    "0000000000", -- linea 674 / direccion 0x2A1 (673) (NOP)
    "0000000000", -- linea 675 / direccion 0x2A2 (674) (NOP)
    "0000000000", -- linea 676 / direccion 0x2A3 (675) (NOP)
    "0000000000", -- linea 677 / direccion 0x2A4 (676) (NOP)
    "0000000000", -- linea 678 / direccion 0x2A5 (677) (NOP)
    "0000000000", -- linea 679 / direccion 0x2A6 (678) (NOP)
    "0000000000", -- linea 680 / direccion 0x2A7 (679) (NOP)
    "0000000000", -- linea 681 / direccion 0x2A8 (680) (NOP)
    "0000000000", -- linea 682 / direccion 0x2A9 (681) (NOP)
    "0000000000", -- linea 683 / direccion 0x2AA (682) (NOP)
    "0000000000", -- linea 684 / direccion 0x2AB (683) (NOP)
    "0000000000", -- linea 685 / direccion 0x2AC (684) (NOP)
    "0000000000", -- linea 686 / direccion 0x2AD (685) (NOP)
    "0000000000", -- linea 687 / direccion 0x2AE (686) (NOP)
    "0000000000", -- linea 688 / direccion 0x2AF (687) (NOP)
    "0000000000", -- linea 689 / direccion 0x2B0 (688) (NOP)
    "0000000000", -- linea 690 / direccion 0x2B1 (689) (NOP)
    "0000000000", -- linea 691 / direccion 0x2B2 (690) (NOP)
    "0000000000", -- linea 692 / direccion 0x2B3 (691) (NOP)
    "0000000000", -- linea 693 / direccion 0x2B4 (692) (NOP)
    "0000000000", -- linea 694 / direccion 0x2B5 (693) (NOP)
    "0000000000", -- linea 695 / direccion 0x2B6 (694) (NOP)
    "0000000000", -- linea 696 / direccion 0x2B7 (695) (NOP)
    "0000000000", -- linea 697 / direccion 0x2B8 (696) (NOP)
    "0000000000", -- linea 698 / direccion 0x2B9 (697) (NOP)
    "0000000000", -- linea 699 / direccion 0x2BA (698) (NOP)
    "0000000000", -- linea 700 / direccion 0x2BB (699) (NOP)
    "0000000000", -- linea 701 / direccion 0x2BC (700) (NOP)
    "0000000000", -- linea 702 / direccion 0x2BD (701) (NOP)
    "0000000000", -- linea 703 / direccion 0x2BE (702) (NOP)
    "0000000000", -- linea 704 / direccion 0x2BF (703) (NOP)
    "0000000000", -- linea 705 / direccion 0x2C0 (704) (NOP)
    "0000000000", -- linea 706 / direccion 0x2C1 (705) (NOP)
    "0000000000", -- linea 707 / direccion 0x2C2 (706) (NOP)
    "0000000000", -- linea 708 / direccion 0x2C3 (707) (NOP)
    "0000000000", -- linea 709 / direccion 0x2C4 (708) (NOP)
    "0000000000", -- linea 710 / direccion 0x2C5 (709) (NOP)
    "0000000000", -- linea 711 / direccion 0x2C6 (710) (NOP)
    "0000000000", -- linea 712 / direccion 0x2C7 (711) (NOP)
    "0000000000", -- linea 713 / direccion 0x2C8 (712) (NOP)
    "0000000000", -- linea 714 / direccion 0x2C9 (713) (NOP)
    "0000000000", -- linea 715 / direccion 0x2CA (714) (NOP)
    "0000000000", -- linea 716 / direccion 0x2CB (715) (NOP)
    "0000000000", -- linea 717 / direccion 0x2CC (716) (NOP)
    "0000000000", -- linea 718 / direccion 0x2CD (717) (NOP)
    "0000000000", -- linea 719 / direccion 0x2CE (718) (NOP)
    "0000000000", -- linea 720 / direccion 0x2CF (719) (NOP)
    "0000000000", -- linea 721 / direccion 0x2D0 (720) (NOP)
    "0000000000", -- linea 722 / direccion 0x2D1 (721) (NOP)
    "0000000000", -- linea 723 / direccion 0x2D2 (722) (NOP)
    "0000000000", -- linea 724 / direccion 0x2D3 (723) (NOP)
    "0000000000", -- linea 725 / direccion 0x2D4 (724) (NOP)
    "0000000000", -- linea 726 / direccion 0x2D5 (725) (NOP)
    "0000000000", -- linea 727 / direccion 0x2D6 (726) (NOP)
    "0000000000", -- linea 728 / direccion 0x2D7 (727) (NOP)
    "0000000000", -- linea 729 / direccion 0x2D8 (728) (NOP)
    "0000000000", -- linea 730 / direccion 0x2D9 (729) (NOP)
    "0000000000", -- linea 731 / direccion 0x2DA (730) (NOP)
    "0000000000", -- linea 732 / direccion 0x2DB (731) (NOP)
    "0000000000", -- linea 733 / direccion 0x2DC (732) (NOP)
    "0000000000", -- linea 734 / direccion 0x2DD (733) (NOP)
    "0000000000", -- linea 735 / direccion 0x2DE (734) (NOP)
    "0000000000", -- linea 736 / direccion 0x2DF (735) (NOP)
    "0000000000", -- linea 737 / direccion 0x2E0 (736) (NOP)
    "0000000000", -- linea 738 / direccion 0x2E1 (737) (NOP)
    "0000000000", -- linea 739 / direccion 0x2E2 (738) (NOP)
    "0000000000", -- linea 740 / direccion 0x2E3 (739) (NOP)
    "0000000000", -- linea 741 / direccion 0x2E4 (740) (NOP)
    "0000000000", -- linea 742 / direccion 0x2E5 (741) (NOP)
    "0000000000", -- linea 743 / direccion 0x2E6 (742) (NOP)
    "0000000000", -- linea 744 / direccion 0x2E7 (743) (NOP)
    "0000000000", -- linea 745 / direccion 0x2E8 (744) (NOP)
    "0000000000", -- linea 746 / direccion 0x2E9 (745) (NOP)
    "0000000000", -- linea 747 / direccion 0x2EA (746) (NOP)
    "0000000000", -- linea 748 / direccion 0x2EB (747) (NOP)
    "0000000000", -- linea 749 / direccion 0x2EC (748) (NOP)
    "0000000000", -- linea 750 / direccion 0x2ED (749) (NOP)
    "0000000000", -- linea 751 / direccion 0x2EE (750) (NOP)
    "0000000000", -- linea 752 / direccion 0x2EF (751) (NOP)
    "0000000000", -- linea 753 / direccion 0x2F0 (752) (NOP)
    "0000000000", -- linea 754 / direccion 0x2F1 (753) (NOP)
    "0000000000", -- linea 755 / direccion 0x2F2 (754) (NOP)
    "0000000000", -- linea 756 / direccion 0x2F3 (755) (NOP)
    "0000000000", -- linea 757 / direccion 0x2F4 (756) (NOP)
    "0000000000", -- linea 758 / direccion 0x2F5 (757) (NOP)
    "0000000000", -- linea 759 / direccion 0x2F6 (758) (NOP)
    "0000000000", -- linea 760 / direccion 0x2F7 (759) (NOP)
    "0000000000", -- linea 761 / direccion 0x2F8 (760) (NOP)
    "0000000000", -- linea 762 / direccion 0x2F9 (761) (NOP)
    "0000000000", -- linea 763 / direccion 0x2FA (762) (NOP)
    "0000000000", -- linea 764 / direccion 0x2FB (763) (NOP)
    "0000000000", -- linea 765 / direccion 0x2FC (764) (NOP)
    "0000000000", -- linea 766 / direccion 0x2FD (765) (NOP)
    "0000000000", -- linea 767 / direccion 0x2FE (766) (NOP)
    "0000000000", -- linea 768 / direccion 0x2FF (767) (NOP)
    "0000000000", -- linea 769 / direccion 0x300 (768) (NOP)
    "0000000000", -- linea 770 / direccion 0x301 (769) (NOP)
    "0000000000", -- linea 771 / direccion 0x302 (770) (NOP)
    "0000000000", -- linea 772 / direccion 0x303 (771) (NOP)
    "0000000000", -- linea 773 / direccion 0x304 (772) (NOP)
    "0000000000", -- linea 774 / direccion 0x305 (773) (NOP)
    "0000000000", -- linea 775 / direccion 0x306 (774) (NOP)
    "0000000000", -- linea 776 / direccion 0x307 (775) (NOP)
    "0000000000", -- linea 777 / direccion 0x308 (776) (NOP)
    "0000000000", -- linea 778 / direccion 0x309 (777) (NOP)
    "0000000000", -- linea 779 / direccion 0x30A (778) (NOP)
    "0000000000", -- linea 780 / direccion 0x30B (779) (NOP)
    "0000000000", -- linea 781 / direccion 0x30C (780) (NOP)
    "0000000000", -- linea 782 / direccion 0x30D (781) (NOP)
    "0000000000", -- linea 783 / direccion 0x30E (782) (NOP)
    "0000000000", -- linea 784 / direccion 0x30F (783) (NOP)
    "0000000000", -- linea 785 / direccion 0x310 (784) (NOP)
    "0000000000", -- linea 786 / direccion 0x311 (785) (NOP)
    "0000000000", -- linea 787 / direccion 0x312 (786) (NOP)
    "0000000000", -- linea 788 / direccion 0x313 (787) (NOP)
    "0000000000", -- linea 789 / direccion 0x314 (788) (NOP)
    "0000000000", -- linea 790 / direccion 0x315 (789) (NOP)
    "0000000000", -- linea 791 / direccion 0x316 (790) (NOP)
    "0000000000", -- linea 792 / direccion 0x317 (791) (NOP)
    "0000000000", -- linea 793 / direccion 0x318 (792) (NOP)
    "0000000000", -- linea 794 / direccion 0x319 (793) (NOP)
    "0000000000", -- linea 795 / direccion 0x31A (794) (NOP)
    "0000000000", -- linea 796 / direccion 0x31B (795) (NOP)
    "0000000000", -- linea 797 / direccion 0x31C (796) (NOP)
    "0000000000", -- linea 798 / direccion 0x31D (797) (NOP)
    "0000000000", -- linea 799 / direccion 0x31E (798) (NOP)
    "0000000000", -- linea 800 / direccion 0x31F (799) (NOP)
    "0000000000", -- linea 801 / direccion 0x320 (800) (NOP)
    "0000000000", -- linea 802 / direccion 0x321 (801) (NOP)
    "0000000000", -- linea 803 / direccion 0x322 (802) (NOP)
    "0000000000", -- linea 804 / direccion 0x323 (803) (NOP)
    "0000000000", -- linea 805 / direccion 0x324 (804) (NOP)
    "0000000000", -- linea 806 / direccion 0x325 (805) (NOP)
    "0000000000", -- linea 807 / direccion 0x326 (806) (NOP)
    "0000000000", -- linea 808 / direccion 0x327 (807) (NOP)
    "0000000000", -- linea 809 / direccion 0x328 (808) (NOP)
    "0000000000", -- linea 810 / direccion 0x329 (809) (NOP)
    "0000000000", -- linea 811 / direccion 0x32A (810) (NOP)
    "0000000000", -- linea 812 / direccion 0x32B (811) (NOP)
    "0000000000", -- linea 813 / direccion 0x32C (812) (NOP)
    "0000000000", -- linea 814 / direccion 0x32D (813) (NOP)
    "0000000000", -- linea 815 / direccion 0x32E (814) (NOP)
    "0000000000", -- linea 816 / direccion 0x32F (815) (NOP)
    "0000000000", -- linea 817 / direccion 0x330 (816) (NOP)
    "0000000000", -- linea 818 / direccion 0x331 (817) (NOP)
    "0000000000", -- linea 819 / direccion 0x332 (818) (NOP)
    "0000000000", -- linea 820 / direccion 0x333 (819) (NOP)
    "0000000000", -- linea 821 / direccion 0x334 (820) (NOP)
    "0000000000", -- linea 822 / direccion 0x335 (821) (NOP)
    "0000000000", -- linea 823 / direccion 0x336 (822) (NOP)
    "0000000000", -- linea 824 / direccion 0x337 (823) (NOP)
    "0000000000", -- linea 825 / direccion 0x338 (824) (NOP)
    "0000000000", -- linea 826 / direccion 0x339 (825) (NOP)
    "0000000000", -- linea 827 / direccion 0x33A (826) (NOP)
    "0000000000", -- linea 828 / direccion 0x33B (827) (NOP)
    "0000000000", -- linea 829 / direccion 0x33C (828) (NOP)
    "0000000000", -- linea 830 / direccion 0x33D (829) (NOP)
    "0000000000", -- linea 831 / direccion 0x33E (830) (NOP)
    "0000000000", -- linea 832 / direccion 0x33F (831) (NOP)
    "0000000000", -- linea 833 / direccion 0x340 (832) (NOP)
    "0000000000", -- linea 834 / direccion 0x341 (833) (NOP)
    "0000000000", -- linea 835 / direccion 0x342 (834) (NOP)
    "0000000000", -- linea 836 / direccion 0x343 (835) (NOP)
    "0000000000", -- linea 837 / direccion 0x344 (836) (NOP)
    "0000000000", -- linea 838 / direccion 0x345 (837) (NOP)
    "0000000000", -- linea 839 / direccion 0x346 (838) (NOP)
    "0000000000", -- linea 840 / direccion 0x347 (839) (NOP)
    "0000000000", -- linea 841 / direccion 0x348 (840) (NOP)
    "0000000000", -- linea 842 / direccion 0x349 (841) (NOP)
    "0000000000", -- linea 843 / direccion 0x34A (842) (NOP)
    "0000000000", -- linea 844 / direccion 0x34B (843) (NOP)
    "0000000000", -- linea 845 / direccion 0x34C (844) (NOP)
    "0000000000", -- linea 846 / direccion 0x34D (845) (NOP)
    "0000000000", -- linea 847 / direccion 0x34E (846) (NOP)
    "0000000000", -- linea 848 / direccion 0x34F (847) (NOP)
    "0000000000", -- linea 849 / direccion 0x350 (848) (NOP)
    "0000000000", -- linea 850 / direccion 0x351 (849) (NOP)
    "0000000000", -- linea 851 / direccion 0x352 (850) (NOP)
    "0000000000", -- linea 852 / direccion 0x353 (851) (NOP)
    "0000000000", -- linea 853 / direccion 0x354 (852) (NOP)
    "0000000000", -- linea 854 / direccion 0x355 (853) (NOP)
    "0000000000", -- linea 855 / direccion 0x356 (854) (NOP)
    "0000000000", -- linea 856 / direccion 0x357 (855) (NOP)
    "0000000000", -- linea 857 / direccion 0x358 (856) (NOP)
    "0000000000", -- linea 858 / direccion 0x359 (857) (NOP)
    "0000000000", -- linea 859 / direccion 0x35A (858) (NOP)
    "0000000000", -- linea 860 / direccion 0x35B (859) (NOP)
    "0000000000", -- linea 861 / direccion 0x35C (860) (NOP)
    "0000000000", -- linea 862 / direccion 0x35D (861) (NOP)
    "0000000000", -- linea 863 / direccion 0x35E (862) (NOP)
    "0000000000", -- linea 864 / direccion 0x35F (863) (NOP)
    "0000000000", -- linea 865 / direccion 0x360 (864) (NOP)
    "0000000000", -- linea 866 / direccion 0x361 (865) (NOP)
    "0000000000", -- linea 867 / direccion 0x362 (866) (NOP)
    "0000000000", -- linea 868 / direccion 0x363 (867) (NOP)
    "0000000000", -- linea 869 / direccion 0x364 (868) (NOP)
    "0000000000", -- linea 870 / direccion 0x365 (869) (NOP)
    "0000000000", -- linea 871 / direccion 0x366 (870) (NOP)
    "0000000000", -- linea 872 / direccion 0x367 (871) (NOP)
    "0000000000", -- linea 873 / direccion 0x368 (872) (NOP)
    "0000000000", -- linea 874 / direccion 0x369 (873) (NOP)
    "0000000000", -- linea 875 / direccion 0x36A (874) (NOP)
    "0000000000", -- linea 876 / direccion 0x36B (875) (NOP)
    "0000000000", -- linea 877 / direccion 0x36C (876) (NOP)
    "0000000000", -- linea 878 / direccion 0x36D (877) (NOP)
    "0000000000", -- linea 879 / direccion 0x36E (878) (NOP)
    "0000000000", -- linea 880 / direccion 0x36F (879) (NOP)
    "0000000000", -- linea 881 / direccion 0x370 (880) (NOP)
    "0000000000", -- linea 882 / direccion 0x371 (881) (NOP)
    "0000000000", -- linea 883 / direccion 0x372 (882) (NOP)
    "0000000000", -- linea 884 / direccion 0x373 (883) (NOP)
    "0000000000", -- linea 885 / direccion 0x374 (884) (NOP)
    "0000000000", -- linea 886 / direccion 0x375 (885) (NOP)
    "0000000000", -- linea 887 / direccion 0x376 (886) (NOP)
    "0000000000", -- linea 888 / direccion 0x377 (887) (NOP)
    "0000000000", -- linea 889 / direccion 0x378 (888) (NOP)
    "0000000000", -- linea 890 / direccion 0x379 (889) (NOP)
    "0000000000", -- linea 891 / direccion 0x37A (890) (NOP)
    "0000000000", -- linea 892 / direccion 0x37B (891) (NOP)
    "0000000000", -- linea 893 / direccion 0x37C (892) (NOP)
    "0000000000", -- linea 894 / direccion 0x37D (893) (NOP)
    "0000000000", -- linea 895 / direccion 0x37E (894) (NOP)
    "0000000000", -- linea 896 / direccion 0x37F (895) (NOP)
    "0000000000", -- linea 897 / direccion 0x380 (896) (NOP)
    "0000000000", -- linea 898 / direccion 0x381 (897) (NOP)
    "0000000000", -- linea 899 / direccion 0x382 (898) (NOP)
    "0000000000", -- linea 900 / direccion 0x383 (899) (NOP)
    "0000000000", -- linea 901 / direccion 0x384 (900) (NOP)
    "0000000000", -- linea 902 / direccion 0x385 (901) (NOP)
    "0000000000", -- linea 903 / direccion 0x386 (902) (NOP)
    "0000000000", -- linea 904 / direccion 0x387 (903) (NOP)
    "0000000000", -- linea 905 / direccion 0x388 (904) (NOP)
    "0000000000", -- linea 906 / direccion 0x389 (905) (NOP)
    "0000000000", -- linea 907 / direccion 0x38A (906) (NOP)
    "0000000000", -- linea 908 / direccion 0x38B (907) (NOP)
    "0000000000", -- linea 909 / direccion 0x38C (908) (NOP)
    "0000000000", -- linea 910 / direccion 0x38D (909) (NOP)
    "0000000000", -- linea 911 / direccion 0x38E (910) (NOP)
    "0000000000", -- linea 912 / direccion 0x38F (911) (NOP)
    "0000000000", -- linea 913 / direccion 0x390 (912) (NOP)
    "0000000000", -- linea 914 / direccion 0x391 (913) (NOP)
    "0000000000", -- linea 915 / direccion 0x392 (914) (NOP)
    "0000000000", -- linea 916 / direccion 0x393 (915) (NOP)
    "0000000000", -- linea 917 / direccion 0x394 (916) (NOP)
    "0000000000", -- linea 918 / direccion 0x395 (917) (NOP)
    "0000000000", -- linea 919 / direccion 0x396 (918) (NOP)
    "0000000000", -- linea 920 / direccion 0x397 (919) (NOP)
    "0000000000", -- linea 921 / direccion 0x398 (920) (NOP)
    "0000000000", -- linea 922 / direccion 0x399 (921) (NOP)
    "0000000000", -- linea 923 / direccion 0x39A (922) (NOP)
    "0000000000", -- linea 924 / direccion 0x39B (923) (NOP)
    "0000000000", -- linea 925 / direccion 0x39C (924) (NOP)
    "0000000000", -- linea 926 / direccion 0x39D (925) (NOP)
    "0000000000", -- linea 927 / direccion 0x39E (926) (NOP)
    "0000000000", -- linea 928 / direccion 0x39F (927) (NOP)
    "0000000000", -- linea 929 / direccion 0x3A0 (928) (NOP)
    "0000000000", -- linea 930 / direccion 0x3A1 (929) (NOP)
    "0000000000", -- linea 931 / direccion 0x3A2 (930) (NOP)
    "0000000000", -- linea 932 / direccion 0x3A3 (931) (NOP)
    "0000000000", -- linea 933 / direccion 0x3A4 (932) (NOP)
    "0000000000", -- linea 934 / direccion 0x3A5 (933) (NOP)
    "0000000000", -- linea 935 / direccion 0x3A6 (934) (NOP)
    "0000000000", -- linea 936 / direccion 0x3A7 (935) (NOP)
    "0000000000", -- linea 937 / direccion 0x3A8 (936) (NOP)
    "0000000000", -- linea 938 / direccion 0x3A9 (937) (NOP)
    "0000000000", -- linea 939 / direccion 0x3AA (938) (NOP)
    "0000000000", -- linea 940 / direccion 0x3AB (939) (NOP)
    "0000000000", -- linea 941 / direccion 0x3AC (940) (NOP)
    "0000000000", -- linea 942 / direccion 0x3AD (941) (NOP)
    "0000000000", -- linea 943 / direccion 0x3AE (942) (NOP)
    "0000000000", -- linea 944 / direccion 0x3AF (943) (NOP)
    "0000000000", -- linea 945 / direccion 0x3B0 (944) (NOP)
    "0000000000", -- linea 946 / direccion 0x3B1 (945) (NOP)
    "0000000000", -- linea 947 / direccion 0x3B2 (946) (NOP)
    "0000000000", -- linea 948 / direccion 0x3B3 (947) (NOP)
    "0000000000", -- linea 949 / direccion 0x3B4 (948) (NOP)
    "0000000000", -- linea 950 / direccion 0x3B5 (949) (NOP)
    "0000000000", -- linea 951 / direccion 0x3B6 (950) (NOP)
    "0000000000", -- linea 952 / direccion 0x3B7 (951) (NOP)
    "0000000000", -- linea 953 / direccion 0x3B8 (952) (NOP)
    "0000000000", -- linea 954 / direccion 0x3B9 (953) (NOP)
    "0000000000", -- linea 955 / direccion 0x3BA (954) (NOP)
    "0000000000", -- linea 956 / direccion 0x3BB (955) (NOP)
    "0000000000", -- linea 957 / direccion 0x3BC (956) (NOP)
    "0000000000", -- linea 958 / direccion 0x3BD (957) (NOP)
    "0000000000", -- linea 959 / direccion 0x3BE (958) (NOP)
    "0000000000", -- linea 960 / direccion 0x3BF (959) (NOP)
    "0000000000", -- linea 961 / direccion 0x3C0 (960) (NOP)
    "0000000000", -- linea 962 / direccion 0x3C1 (961) (NOP)
    "0000000000", -- linea 963 / direccion 0x3C2 (962) (NOP)
    "0000000000", -- linea 964 / direccion 0x3C3 (963) (NOP)
    "0000000000", -- linea 965 / direccion 0x3C4 (964) (NOP)
    "0000000000", -- linea 966 / direccion 0x3C5 (965) (NOP)
    "0000000000", -- linea 967 / direccion 0x3C6 (966) (NOP)
    "0000000000", -- linea 968 / direccion 0x3C7 (967) (NOP)
    "0000000000", -- linea 969 / direccion 0x3C8 (968) (NOP)
    "0000000000", -- linea 970 / direccion 0x3C9 (969) (NOP)
    "0000000000", -- linea 971 / direccion 0x3CA (970) (NOP)
    "0000000000", -- linea 972 / direccion 0x3CB (971) (NOP)
    "0000000000", -- linea 973 / direccion 0x3CC (972) (NOP)
    "0000000000", -- linea 974 / direccion 0x3CD (973) (NOP)
    "0000000000", -- linea 975 / direccion 0x3CE (974) (NOP)
    "0000000000", -- linea 976 / direccion 0x3CF (975) (NOP)
    "0000000000", -- linea 977 / direccion 0x3D0 (976) (NOP)
    "0000000000", -- linea 978 / direccion 0x3D1 (977) (NOP)
    "0000000000", -- linea 979 / direccion 0x3D2 (978) (NOP)
    "0000000000", -- linea 980 / direccion 0x3D3 (979) (NOP)
    "0000000000", -- linea 981 / direccion 0x3D4 (980) (NOP)
    "0000000000", -- linea 982 / direccion 0x3D5 (981) (NOP)
    "0000000000", -- linea 983 / direccion 0x3D6 (982) (NOP)
    "0000000000", -- linea 984 / direccion 0x3D7 (983) (NOP)
    "0000000000", -- linea 985 / direccion 0x3D8 (984) (NOP)
    "0000000000", -- linea 986 / direccion 0x3D9 (985) (NOP)
    "0000000000", -- linea 987 / direccion 0x3DA (986) (NOP)
    "0000000000", -- linea 988 / direccion 0x3DB (987) (NOP)
    "0000000000", -- linea 989 / direccion 0x3DC (988) (NOP)
    "0000000000", -- linea 990 / direccion 0x3DD (989) (NOP)
    "0000000000", -- linea 991 / direccion 0x3DE (990) (NOP)
    "0000000000", -- linea 992 / direccion 0x3DF (991) (NOP)
    "0000000000", -- linea 993 / direccion 0x3E0 (992) (NOP)
    "0000000000", -- linea 994 / direccion 0x3E1 (993) (NOP)
    "0000000000", -- linea 995 / direccion 0x3E2 (994) (NOP)
    "0000000000", -- linea 996 / direccion 0x3E3 (995) (NOP)
    "0000000000", -- linea 997 / direccion 0x3E4 (996) (NOP)
    "0000000000", -- linea 998 / direccion 0x3E5 (997) (NOP)
    "0000000000", -- linea 999 / direccion 0x3E6 (998) (NOP)
    "0000000000", -- linea 1000 / direccion 0x3E7 (999) (NOP)
    "0000000000", -- linea 1001 / direccion 0x3E8 (1000) (NOP)
    "0000000000", -- linea 1002 / direccion 0x3E9 (1001) (NOP)
    "0000000000", -- linea 1003 / direccion 0x3EA (1002) (NOP)
    "0000000000", -- linea 1004 / direccion 0x3EB (1003) (NOP)
    "0000000000", -- linea 1005 / direccion 0x3EC (1004) (NOP)
    "0000000000", -- linea 1006 / direccion 0x3ED (1005) (NOP)
    "0000000000", -- linea 1007 / direccion 0x3EE (1006) (NOP)
    "0000000000", -- linea 1008 / direccion 0x3EF (1007) (NOP)
    "0000000000", -- linea 1009 / direccion 0x3F0 (1008) (NOP)
    "0000000000", -- linea 1010 / direccion 0x3F1 (1009) (NOP)
    "0000000000", -- linea 1011 / direccion 0x3F2 (1010) (NOP)
    "0000000000", -- linea 1012 / direccion 0x3F3 (1011) (NOP)
    "0000000000", -- linea 1013 / direccion 0x3F4 (1012) (NOP)
    "0000000000", -- linea 1014 / direccion 0x3F5 (1013) (NOP)
    "0000000000", -- linea 1015 / direccion 0x3F6 (1014) (NOP)
    "0000000000", -- linea 1016 / direccion 0x3F7 (1015) (NOP)
    "0000000000", -- linea 1017 / direccion 0x3F8 (1016) (NOP)
    "0000000000", -- linea 1018 / direccion 0x3F9 (1017) (NOP)
    "0000000000", -- linea 1019 / direccion 0x3FA (1018) (NOP)
    "0000000000", -- linea 1020 / direccion 0x3FB (1019) (NOP)
    "0000000000", -- linea 1021 / direccion 0x3FC (1020) (NOP)
    "0000000000", -- linea 1022 / direccion 0x3FD (1021) (NOP)
    "0000000000", -- linea 1023 / direccion 0x3FE (1022) (NOP)
    "0000000000", -- linea 1024 / direccion 0x3FF (1023) (NOP)
	others => (others => '0')
	);

begin

	data <= ROM(to_integer(unsigned(addr)));

end arq1;
