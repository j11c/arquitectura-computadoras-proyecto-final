-------------------------------------------------------------------------------
--
-- Company : Universidad Miguel Hernandez
-- Engineer: joshi
-- 
-- Create Date:    20/11/2025 13:45:11
-- Project Name:   UnidadControl
-- Module Name:    UnidadControl.vhd
-- Description:
--
-- Additional Comments:
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;  -- Para std_logic
use IEEE.numeric_std.all;     -- Para unsigned

entity UnidadControl is
	port(
		clk 	: in std_logic;
		instr 	: in std_logic_vector(9 downto 0);
		ctrl 	: out std_logic_vector(12 downto 0)
	);
end UnidadControl;

architecture arq1 of UnidadControl is

	-- Estructuras de memorias
	type memOper2Param is array(0 to 512) of std_logic_vector(15 downto 0);
	type memOper1Param is array(0 to 512) of std_logic_vector(15 downto 0);
	type memIndirecto is array(0 to 512) of std_logic_vector(15 downto 0);

	-- Contenidos
	signal Oper2Param : memOper2Param := (
		-- MODO 00
		x"0100", x"0280", x"1008", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER A, A
		x"0100", x"0280", x"1008", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER A, B
		x"0100", x"0280", x"1008", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER A, C
		x"0100", x"0280", x"1008", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER A, D
		x"0100", x"0280", x"1004", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER B, A
		x"0100", x"0280", x"1004", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER B, B
		x"0100", x"0280", x"1004", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER B, C
		x"0100", x"0280", x"1004", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER B, D
		x"0100", x"0280", x"1002", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER C, A
		x"0100", x"0280", x"1002", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER C, B
		x"0100", x"0280", x"1002", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER C, C
		x"0100", x"0280", x"1002", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER C, D
		x"0100", x"0280", x"1001", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER D, A
		x"0100", x"0280", x"1001", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER D, B
		x"0100", x"0280", x"1001", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER D, C
		x"0100", x"0280", x"1001", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER D, D
		-- MODO 01
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1008", x"0000", x"0000", -- OPER A, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1008", x"0000", x"0000", -- OPER A, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1008", x"0000", x"0000", -- OPER A, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1008", x"0000", x"0000", -- OPER A, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1004", x"0000", x"0000", -- OPER B, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1004", x"0000", x"0000", -- OPER B, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1004", x"0000", x"0000", -- OPER B, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1004", x"0000", x"0000", -- OPER B, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1002", x"0000", x"0000", -- OPER C, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1002", x"0000", x"0000", -- OPER C, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1002", x"0000", x"0000", -- OPER C, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1002", x"0000", x"0000", -- OPER C, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1001", x"0000", x"0000", -- OPER D, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1001", x"0000", x"0000", -- OPER D, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1001", x"0000", x"0000", -- OPER D, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1001", x"0000", x"0000", -- OPER D, [DIR]
		-- MODO 10
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR], A
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR], A
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR], A
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR], A
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR], B
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR], B
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR], B
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR], B
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR], C
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR], C
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR], C
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR], C
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR], D
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR], D
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR], D
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR], D
		-- MODO 11
		x"0100", x"0280", x"0100", x"0240", x"1008", x"0000", x"0000", x"0000", -- OPER A, #num
		x"0100", x"0280", x"0100", x"0240", x"1008", x"0000", x"0000", x"0000", -- OPER A, #num
		x"0100", x"0280", x"0100", x"0240", x"1008", x"0000", x"0000", x"0000", -- OPER A, #num
		x"0100", x"0280", x"0100", x"0240", x"1008", x"0000", x"0000", x"0000", -- OPER A, #num
		x"0100", x"0280", x"0100", x"0240", x"1004", x"0000", x"0000", x"0000", -- OPER B, #num
		x"0100", x"0280", x"0100", x"0240", x"1004", x"0000", x"0000", x"0000", -- OPER B, #num
		x"0100", x"0280", x"0100", x"0240", x"1004", x"0000", x"0000", x"0000", -- OPER B, #num
		x"0100", x"0280", x"0100", x"0240", x"1004", x"0000", x"0000", x"0000", -- OPER B, #num
		x"0100", x"0280", x"0100", x"0240", x"1002", x"0000", x"0000", x"0000", -- OPER C, #num
		x"0100", x"0280", x"0100", x"0240", x"1002", x"0000", x"0000", x"0000", -- OPER C, #num
		x"0100", x"0280", x"0100", x"0240", x"1002", x"0000", x"0000", x"0000", -- OPER C, #num
		x"0100", x"0280", x"0100", x"0240", x"1002", x"0000", x"0000", x"0000", -- OPER C, #num
		x"0100", x"0280", x"0100", x"0240", x"1001", x"0000", x"0000", x"0000", -- OPER D, #num
		x"0100", x"0280", x"0100", x"0240", x"1001", x"0000", x"0000", x"0000", -- OPER D, #num
		x"0100", x"0280", x"0100", x"0240", x"1001", x"0000", x"0000", x"0000", -- OPER D, #num
		x"0100", x"0280", x"0100", x"0240", x"1001", x"0000", x"0000", x"0000", -- OPER D, #num
		others => x"00000"
	);
	
	signal Comparacion : memOper2Param := (
		-- MODO 00
		x"0100", x"0280", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER A, A
		x"0100", x"0280", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER A, B
		x"0100", x"0280", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER A, C
		x"0100", x"0280", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER A, D
		x"0100", x"0280", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER B, A
		x"0100", x"0280", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER B, B
		x"0100", x"0280", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER B, C
		x"0100", x"0280", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER B, D
		x"0100", x"0280", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER C, A
		x"0100", x"0280", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER C, B
		x"0100", x"0280", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER C, C
		x"0100", x"0280", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER C, D
		x"0100", x"0280", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER D, A
		x"0100", x"0280", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER D, B
		x"0100", x"0280", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER D, C
		x"0100", x"0280", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER D, D
		-- MODO 01
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER A, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER A, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER A, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER A, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER B, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER B, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER B, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER B, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER C, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER C, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER C, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER C, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER D, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER D, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER D, [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER D, [DIR]
		-- MODO 10
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER [DIR], A
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER [DIR], A
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER [DIR], A
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER [DIR], A
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER [DIR], B
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER [DIR], B
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER [DIR], B
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER [DIR], B
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER [DIR], C
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER [DIR], C
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER [DIR], C
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER [DIR], C
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER [DIR], D
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER [DIR], D
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER [DIR], D
		x"0100", x"0280", x"0100", x"0220", x"0040", x"0000", x"0000", x"0000", -- OPER [DIR], D
		-- MODO 11
		x"0100", x"0280", x"0100", x"0240", x"0000", x"0000", x"0000", x"0000", -- OPER A, #num
		x"0100", x"0280", x"0100", x"0240", x"0000", x"0000", x"0000", x"0000", -- OPER A, #num
		x"0100", x"0280", x"0100", x"0240", x"0000", x"0000", x"0000", x"0000", -- OPER A, #num
		x"0100", x"0280", x"0100", x"0240", x"0000", x"0000", x"0000", x"0000", -- OPER A, #num
		x"0100", x"0280", x"0100", x"0240", x"0000", x"0000", x"0000", x"0000", -- OPER B, #num
		x"0100", x"0280", x"0100", x"0240", x"0000", x"0000", x"0000", x"0000", -- OPER B, #num
		x"0100", x"0280", x"0100", x"0240", x"0000", x"0000", x"0000", x"0000", -- OPER B, #num
		x"0100", x"0280", x"0100", x"0240", x"0000", x"0000", x"0000", x"0000", -- OPER B, #num
		x"0100", x"0280", x"0100", x"0240", x"0000", x"0000", x"0000", x"0000", -- OPER C, #num
		x"0100", x"0280", x"0100", x"0240", x"0000", x"0000", x"0000", x"0000", -- OPER C, #num
		x"0100", x"0280", x"0100", x"0240", x"0000", x"0000", x"0000", x"0000", -- OPER C, #num
		x"0100", x"0280", x"0100", x"0240", x"0000", x"0000", x"0000", x"0000", -- OPER C, #num
		x"0100", x"0280", x"0100", x"0240", x"0000", x"0000", x"0000", x"0000", -- OPER D, #num
		x"0100", x"0280", x"0100", x"0240", x"0000", x"0000", x"0000", x"0000", -- OPER D, #num
		x"0100", x"0280", x"0100", x"0240", x"0000", x"0000", x"0000", x"0000", -- OPER D, #num
		x"0100", x"0280", x"0100", x"0240", x"0000", x"0000", x"0000", x"0000", -- OPER D, #num
		others => x"00000"
	);

	signal Oper1Param : memOper1Param := (
		-- MODO 00
		x"0100", x"0280", x"1008", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER A
		x"0100", x"0280", x"1004", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER B
		x"0100", x"0280", x"1002", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER C
		x"0100", x"0280", x"1001", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER D
		x"0100", x"0280", x"1008", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER A
		x"0100", x"0280", x"1004", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER B
		x"0100", x"0280", x"1002", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER C
		x"0100", x"0280", x"1001", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER D
		x"0100", x"0280", x"1008", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER A
		x"0100", x"0280", x"1004", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER B
		x"0100", x"0280", x"1002", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER C
		x"0100", x"0280", x"1001", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER D
		x"0100", x"0280", x"1008", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER A
		x"0100", x"0280", x"1004", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER B
		x"0100", x"0280", x"1002", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER C
		x"0100", x"0280", x"1001", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER D

		-- MODO 01
		x"0100", x"0280", x"1008", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER A
		x"0100", x"0280", x"1004", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER B
		x"0100", x"0280", x"1002", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER C
		x"0100", x"0280", x"1001", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER D
		x"0100", x"0280", x"1008", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER A
		x"0100", x"0280", x"1004", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER B
		x"0100", x"0280", x"1002", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER C
		x"0100", x"0280", x"1001", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER D
		x"0100", x"0280", x"1008", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER A
		x"0100", x"0280", x"1004", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER B
		x"0100", x"0280", x"1002", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER C
		x"0100", x"0280", x"1001", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER D
		x"0100", x"0280", x"1008", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER A
		x"0100", x"0280", x"1004", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER B
		x"0100", x"0280", x"1002", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER C
		x"0100", x"0280", x"1001", x"0000", x"0000", x"0000", x"0000", x"0000", -- OPER D

		-- MODO 10 (memoria)
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]

		-- MODO 11 (memoria)
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		x"0100", x"0280", x"0100", x"0220", x"0040", x"1010", x"0000", x"0000", -- OPER [DIR]
		others => x"00000"
	);

	signal Saltos 	  : memOper2Param := (
		-- MODO 00 JMP
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JMP [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JMP [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JMP [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JMP [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JMP [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JMP [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JMP [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JMP [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JMP [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JMP [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JMP [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JMP [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JMP [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JMP [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JMP [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JMP [DIR]

		-- MODO 01 JLT
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JLT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JLT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JLT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JLT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JLT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JLT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JLT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JLT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JLT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JLT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JLT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JLT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JLT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JLT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JLT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JLT [DIR]

		-- MODO 10 JGT
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JGT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JGT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JGT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JGT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JGT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JGT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JGT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JGT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JGT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JGT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JGT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JGT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JGT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JGT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JGT [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JGT [DIR]

		-- MODO 11 JEQ
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JEQ [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JEQ [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JEQ [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JEQ [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JEQ [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JEQ [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JEQ [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JEQ [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JEQ [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JEQ [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JEQ [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JEQ [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JEQ [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JEQ [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JEQ [DIR]
		x"0100", x"0280", x"0100", x"1400", x"0000", x"0000", x"0000", x"0000", -- JEQ [DIR]
		others => x"00000"
	);

	signal Indirecto  : memIndirecto  := (
		-- MODO 00
		x"0100", x"0280", x"0020", x"0040", x"1008", x"0000", x"0000", x"0000", -- ILOAD A, [A]
		x"0100", x"0280", x"0020", x"0040", x"1008", x"0000", x"0000", x"0000", -- ILOAD A, [B]
		x"0100", x"0280", x"0020", x"0040", x"1008", x"0000", x"0000", x"0000", -- ILOAD A, [C]
		x"0100", x"0280", x"0020", x"0040", x"1008", x"0000", x"0000", x"0000", -- ILOAD A, [D]
		x"0100", x"0280", x"0020", x"0040", x"1004", x"0000", x"0000", x"0000", -- ILOAD B, [A]
		x"0100", x"0280", x"0020", x"0040", x"1004", x"0000", x"0000", x"0000", -- ILOAD B, [B]
		x"0100", x"0280", x"0020", x"0040", x"1004", x"0000", x"0000", x"0000", -- ILOAD B, [C]
		x"0100", x"0280", x"0020", x"0040", x"1004", x"0000", x"0000", x"0000", -- ILOAD B, [D]
		x"0100", x"0280", x"0020", x"0040", x"1002", x"0000", x"0000", x"0000", -- ILOAD C, [A]
		x"0100", x"0280", x"0020", x"0040", x"1002", x"0000", x"0000", x"0000", -- ILOAD C, [B]
		x"0100", x"0280", x"0020", x"0040", x"1002", x"0000", x"0000", x"0000", -- ILOAD C, [C]
		x"0100", x"0280", x"0020", x"0040", x"1002", x"0000", x"0000", x"0000", -- ILOAD C, [D]
		x"0100", x"0280", x"0020", x"0040", x"1001", x"0000", x"0000", x"0000", -- ILOAD D, [A]
		x"0100", x"0280", x"0020", x"0040", x"1001", x"0000", x"0000", x"0000", -- ILOAD D, [B]
		x"0100", x"0280", x"0020", x"0040", x"1001", x"0000", x"0000", x"0000", -- ILOAD D, [C]
		x"0100", x"0280", x"0020", x"0040", x"1001", x"0000", x"0000", x"0000", -- ILOAD D, [D]
		others => x"00000"
	);

	-- FALTA ENTRADA Y SALIDA

	signal control_signals : std_logic_vector(15 downto 0) := (others => '0');
	signal microCounter : unsigned(2 downto 0) := (others => '0');
	signal addr : std_logic_vector(8 downto 0) := (others => '0');
	signal coop : std_logic_vector(3 downto 0) := (others => '0');
	
begin
	
	coop <= instr(9 downto 6);
	addr <= instr(5 downto 0) & std_logic_vector(microCounter);
	
	with coop select control_signals <= 
		Oper2Param(to_integer(unsigned(addr))) when "0001", -- ADD
		Oper2Param(to_integer(unsigned(addr))) when "0010", -- SUB
		Oper2Param(to_integer(unsigned(addr))) when "0011", -- MUL
		Oper2Param(to_integer(unsigned(addr))) when "0100", -- DIV
		Oper2Param(to_integer(unsigned(addr))) when "0101", -- AND
		Oper2Param(to_integer(unsigned(addr))) when "0110", -- OR
		Oper2Param(to_integer(unsigned(addr))) when "1001", -- LOAD

		Comparacion(to_integer(unsigned(addr))) when "1000", -- CMP

		Oper1Param(to_integer(unsigned(addr))) when "0111", -- NOT
		Oper1Param(to_integer(unsigned(addr))) when "1010", -- INC/DEC
		Oper1Param(to_integer(unsigned(addr))) when "1011", -- SHL/SHR

		Saltos(to_integer(unsigned(addr))) when "1101",

--		Oper1Param(to_integer(unsigned(addr))) when "0000", -- HALT

		Indirecto(to_integer(unsigned(addr))) when "1110",
		x"00000" when others;

	process (clk, Instr, control_signals, addr)
	begin
		ctrl <= control_signals(12 downto 0);
		if rising_edge(clk) then
			microCounter + 1;
		end if;
	end process;

end arq1;
