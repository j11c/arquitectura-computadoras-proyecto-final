-------------------------------------------------------------------------------
--
-- Company : Universidad Miguel Hernandez
-- Engineer: joshi
-- 
-- Create Date:    20/11/2025 09:37:07
-- Project Name:   memoriaPrograma
-- Module Name:    memoriaPrograma.vhd
-- Description:
--
-- Additional Comments:
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;  -- Para std_logic
use IEEE.numeric_std.all;     -- Para unsigned

entity memoriaPrograma is
	port( 
		addr : in  std_logic_vector(9 downto 0);
        data : out std_logic_vector(9 downto 0)
	);
end memoriaPrograma;

architecture arq1 of memoriaPrograma is
	
	type mem_type is array (0 to 1023) of std_logic_vector(9 downto 0);

	constant ROM : mem_type := (
"1001110000", -- linea 1 / direccion 0
"0000000101", -- linea 2 / direccion 1
"1100100000", -- linea 3 / direccion 2
"0000000000", -- linea 4 / direccion 3
"1111000000", -- linea 5 / direccion 4 (NOP)
"1111000000", -- linea 6 / direccion 5 (NOP)
"1111000000", -- linea 7 / direccion 6 (NOP)
"1111000000", -- linea 8 / direccion 7 (NOP)
"1111000000", -- linea 9 / direccion 8 (NOP)
"1111000000", -- linea 10 / direccion 9 (NOP)
"1111000000", -- linea 11 / direccion 10 (NOP)
"1111000000", -- linea 12 / direccion 11 (NOP)
"1111000000", -- linea 13 / direccion 12 (NOP)
"1111000000", -- linea 14 / direccion 13 (NOP)
"1111000000", -- linea 15 / direccion 14 (NOP)
"1111000000", -- linea 16 / direccion 15 (NOP)
"1111000000", -- linea 17 / direccion 16 (NOP)
"1111000000", -- linea 18 / direccion 17 (NOP)
"1111000000", -- linea 19 / direccion 18 (NOP)
"1111000000", -- linea 20 / direccion 19 (NOP)
"1111000000", -- linea 21 / direccion 20 (NOP)
"1111000000", -- linea 22 / direccion 21 (NOP)
"1111000000", -- linea 23 / direccion 22 (NOP)
"1111000000", -- linea 24 / direccion 23 (NOP)
"1111000000", -- linea 25 / direccion 24 (NOP)
"1111000000", -- linea 26 / direccion 25 (NOP)
"1111000000", -- linea 27 / direccion 26 (NOP)
"1111000000", -- linea 28 / direccion 27 (NOP)
"1111000000", -- linea 29 / direccion 28 (NOP)
"1111000000", -- linea 30 / direccion 29 (NOP)
"1111000000", -- linea 31 / direccion 30 (NOP)
"1111000000", -- linea 32 / direccion 31 (NOP)
"1111000000", -- linea 33 / direccion 32 (NOP)
"1111000000", -- linea 34 / direccion 33 (NOP)
"1111000000", -- linea 35 / direccion 34 (NOP)
"1111000000", -- linea 36 / direccion 35 (NOP)
"1111000000", -- linea 37 / direccion 36 (NOP)
"1111000000", -- linea 38 / direccion 37 (NOP)
"1111000000", -- linea 39 / direccion 38 (NOP)
"1111000000", -- linea 40 / direccion 39 (NOP)
"1111000000", -- linea 41 / direccion 40 (NOP)
"1111000000", -- linea 42 / direccion 41 (NOP)
"1111000000", -- linea 43 / direccion 42 (NOP)
"1111000000", -- linea 44 / direccion 43 (NOP)
"1111000000", -- linea 45 / direccion 44 (NOP)
"1111000000", -- linea 46 / direccion 45 (NOP)
"1111000000", -- linea 47 / direccion 46 (NOP)
"1111000000", -- linea 48 / direccion 47 (NOP)
"1111000000", -- linea 49 / direccion 48 (NOP)
"1111000000", -- linea 50 / direccion 49 (NOP)
"1111000000", -- linea 51 / direccion 50 (NOP)
"1111000000", -- linea 52 / direccion 51 (NOP)
"1111000000", -- linea 53 / direccion 52 (NOP)
"1111000000", -- linea 54 / direccion 53 (NOP)
"1111000000", -- linea 55 / direccion 54 (NOP)
"1111000000", -- linea 56 / direccion 55 (NOP)
"1111000000", -- linea 57 / direccion 56 (NOP)
"1111000000", -- linea 58 / direccion 57 (NOP)
"1111000000", -- linea 59 / direccion 58 (NOP)
"1111000000", -- linea 60 / direccion 59 (NOP)
"1111000000", -- linea 61 / direccion 60 (NOP)
"1111000000", -- linea 62 / direccion 61 (NOP)
"1111000000", -- linea 63 / direccion 62 (NOP)
"1111000000", -- linea 64 / direccion 63 (NOP)
"1111000000", -- linea 65 / direccion 64 (NOP)
"1111000000", -- linea 66 / direccion 65 (NOP)
"1111000000", -- linea 67 / direccion 66 (NOP)
"1111000000", -- linea 68 / direccion 67 (NOP)
"1111000000", -- linea 69 / direccion 68 (NOP)
"1111000000", -- linea 70 / direccion 69 (NOP)
"1111000000", -- linea 71 / direccion 70 (NOP)
"1111000000", -- linea 72 / direccion 71 (NOP)
"1111000000", -- linea 73 / direccion 72 (NOP)
"1111000000", -- linea 74 / direccion 73 (NOP)
"1111000000", -- linea 75 / direccion 74 (NOP)
"1111000000", -- linea 76 / direccion 75 (NOP)
"1111000000", -- linea 77 / direccion 76 (NOP)
"1111000000", -- linea 78 / direccion 77 (NOP)
"1111000000", -- linea 79 / direccion 78 (NOP)
"1111000000", -- linea 80 / direccion 79 (NOP)
"1111000000", -- linea 81 / direccion 80 (NOP)
"1111000000", -- linea 82 / direccion 81 (NOP)
"1111000000", -- linea 83 / direccion 82 (NOP)
"1111000000", -- linea 84 / direccion 83 (NOP)
"1111000000", -- linea 85 / direccion 84 (NOP)
"1111000000", -- linea 86 / direccion 85 (NOP)
"1111000000", -- linea 87 / direccion 86 (NOP)
"1111000000", -- linea 88 / direccion 87 (NOP)
"1111000000", -- linea 89 / direccion 88 (NOP)
"1111000000", -- linea 90 / direccion 89 (NOP)
"1111000000", -- linea 91 / direccion 90 (NOP)
"1111000000", -- linea 92 / direccion 91 (NOP)
"1111000000", -- linea 93 / direccion 92 (NOP)
"1111000000", -- linea 94 / direccion 93 (NOP)
"1111000000", -- linea 95 / direccion 94 (NOP)
"1111000000", -- linea 96 / direccion 95 (NOP)
"1111000000", -- linea 97 / direccion 96 (NOP)
"1111000000", -- linea 98 / direccion 97 (NOP)
"1111000000", -- linea 99 / direccion 98 (NOP)
"1111000000", -- linea 100 / direccion 99 (NOP)
"1111000000", -- linea 101 / direccion 100 (NOP)
"1111000000", -- linea 102 / direccion 101 (NOP)
"1111000000", -- linea 103 / direccion 102 (NOP)
"1111000000", -- linea 104 / direccion 103 (NOP)
"1111000000", -- linea 105 / direccion 104 (NOP)
"1111000000", -- linea 106 / direccion 105 (NOP)
"1111000000", -- linea 107 / direccion 106 (NOP)
"1111000000", -- linea 108 / direccion 107 (NOP)
"1111000000", -- linea 109 / direccion 108 (NOP)
"1111000000", -- linea 110 / direccion 109 (NOP)
"1111000000", -- linea 111 / direccion 110 (NOP)
"1111000000", -- linea 112 / direccion 111 (NOP)
"1111000000", -- linea 113 / direccion 112 (NOP)
"1111000000", -- linea 114 / direccion 113 (NOP)
"1111000000", -- linea 115 / direccion 114 (NOP)
"1111000000", -- linea 116 / direccion 115 (NOP)
"1111000000", -- linea 117 / direccion 116 (NOP)
"1111000000", -- linea 118 / direccion 117 (NOP)
"1111000000", -- linea 119 / direccion 118 (NOP)
"1111000000", -- linea 120 / direccion 119 (NOP)
"1111000000", -- linea 121 / direccion 120 (NOP)
"1111000000", -- linea 122 / direccion 121 (NOP)
"1111000000", -- linea 123 / direccion 122 (NOP)
"1111000000", -- linea 124 / direccion 123 (NOP)
"1111000000", -- linea 125 / direccion 124 (NOP)
"1111000000", -- linea 126 / direccion 125 (NOP)
"1111000000", -- linea 127 / direccion 126 (NOP)
"1111000000", -- linea 128 / direccion 127 (NOP)
"1111000000", -- linea 129 / direccion 128 (NOP)
"1111000000", -- linea 130 / direccion 129 (NOP)
"1111000000", -- linea 131 / direccion 130 (NOP)
"1111000000", -- linea 132 / direccion 131 (NOP)
"1111000000", -- linea 133 / direccion 132 (NOP)
"1111000000", -- linea 134 / direccion 133 (NOP)
"1111000000", -- linea 135 / direccion 134 (NOP)
"1111000000", -- linea 136 / direccion 135 (NOP)
"1111000000", -- linea 137 / direccion 136 (NOP)
"1111000000", -- linea 138 / direccion 137 (NOP)
"1111000000", -- linea 139 / direccion 138 (NOP)
"1111000000", -- linea 140 / direccion 139 (NOP)
"1111000000", -- linea 141 / direccion 140 (NOP)
"1111000000", -- linea 142 / direccion 141 (NOP)
"1111000000", -- linea 143 / direccion 142 (NOP)
"1111000000", -- linea 144 / direccion 143 (NOP)
"1111000000", -- linea 145 / direccion 144 (NOP)
"1111000000", -- linea 146 / direccion 145 (NOP)
"1111000000", -- linea 147 / direccion 146 (NOP)
"1111000000", -- linea 148 / direccion 147 (NOP)
"1111000000", -- linea 149 / direccion 148 (NOP)
"1111000000", -- linea 150 / direccion 149 (NOP)
"1111000000", -- linea 151 / direccion 150 (NOP)
"1111000000", -- linea 152 / direccion 151 (NOP)
"1111000000", -- linea 153 / direccion 152 (NOP)
"1111000000", -- linea 154 / direccion 153 (NOP)
"1111000000", -- linea 155 / direccion 154 (NOP)
"1111000000", -- linea 156 / direccion 155 (NOP)
"1111000000", -- linea 157 / direccion 156 (NOP)
"1111000000", -- linea 158 / direccion 157 (NOP)
"1111000000", -- linea 159 / direccion 158 (NOP)
"1111000000", -- linea 160 / direccion 159 (NOP)
"1111000000", -- linea 161 / direccion 160 (NOP)
"1111000000", -- linea 162 / direccion 161 (NOP)
"1111000000", -- linea 163 / direccion 162 (NOP)
"1111000000", -- linea 164 / direccion 163 (NOP)
"1111000000", -- linea 165 / direccion 164 (NOP)
"1111000000", -- linea 166 / direccion 165 (NOP)
"1111000000", -- linea 167 / direccion 166 (NOP)
"1111000000", -- linea 168 / direccion 167 (NOP)
"1111000000", -- linea 169 / direccion 168 (NOP)
"1111000000", -- linea 170 / direccion 169 (NOP)
"1111000000", -- linea 171 / direccion 170 (NOP)
"1111000000", -- linea 172 / direccion 171 (NOP)
"1111000000", -- linea 173 / direccion 172 (NOP)
"1111000000", -- linea 174 / direccion 173 (NOP)
"1111000000", -- linea 175 / direccion 174 (NOP)
"1111000000", -- linea 176 / direccion 175 (NOP)
"1111000000", -- linea 177 / direccion 176 (NOP)
"1111000000", -- linea 178 / direccion 177 (NOP)
"1111000000", -- linea 179 / direccion 178 (NOP)
"1111000000", -- linea 180 / direccion 179 (NOP)
"1111000000", -- linea 181 / direccion 180 (NOP)
"1111000000", -- linea 182 / direccion 181 (NOP)
"1111000000", -- linea 183 / direccion 182 (NOP)
"1111000000", -- linea 184 / direccion 183 (NOP)
"1111000000", -- linea 185 / direccion 184 (NOP)
"1111000000", -- linea 186 / direccion 185 (NOP)
"1111000000", -- linea 187 / direccion 186 (NOP)
"1111000000", -- linea 188 / direccion 187 (NOP)
"1111000000", -- linea 189 / direccion 188 (NOP)
"1111000000", -- linea 190 / direccion 189 (NOP)
"1111000000", -- linea 191 / direccion 190 (NOP)
"1111000000", -- linea 192 / direccion 191 (NOP)
"1111000000", -- linea 193 / direccion 192 (NOP)
"1111000000", -- linea 194 / direccion 193 (NOP)
"1111000000", -- linea 195 / direccion 194 (NOP)
"1111000000", -- linea 196 / direccion 195 (NOP)
"1111000000", -- linea 197 / direccion 196 (NOP)
"1111000000", -- linea 198 / direccion 197 (NOP)
"1111000000", -- linea 199 / direccion 198 (NOP)
"1111000000", -- linea 200 / direccion 199 (NOP)
"1111000000", -- linea 201 / direccion 200 (NOP)
"1111000000", -- linea 202 / direccion 201 (NOP)
"1111000000", -- linea 203 / direccion 202 (NOP)
"1111000000", -- linea 204 / direccion 203 (NOP)
"1111000000", -- linea 205 / direccion 204 (NOP)
"1111000000", -- linea 206 / direccion 205 (NOP)
"1111000000", -- linea 207 / direccion 206 (NOP)
"1111000000", -- linea 208 / direccion 207 (NOP)
"1111000000", -- linea 209 / direccion 208 (NOP)
"1111000000", -- linea 210 / direccion 209 (NOP)
"1111000000", -- linea 211 / direccion 210 (NOP)
"1111000000", -- linea 212 / direccion 211 (NOP)
"1111000000", -- linea 213 / direccion 212 (NOP)
"1111000000", -- linea 214 / direccion 213 (NOP)
"1111000000", -- linea 215 / direccion 214 (NOP)
"1111000000", -- linea 216 / direccion 215 (NOP)
"1111000000", -- linea 217 / direccion 216 (NOP)
"1111000000", -- linea 218 / direccion 217 (NOP)
"1111000000", -- linea 219 / direccion 218 (NOP)
"1111000000", -- linea 220 / direccion 219 (NOP)
"1111000000", -- linea 221 / direccion 220 (NOP)
"1111000000", -- linea 222 / direccion 221 (NOP)
"1111000000", -- linea 223 / direccion 222 (NOP)
"1111000000", -- linea 224 / direccion 223 (NOP)
"1111000000", -- linea 225 / direccion 224 (NOP)
"1111000000", -- linea 226 / direccion 225 (NOP)
"1111000000", -- linea 227 / direccion 226 (NOP)
"1111000000", -- linea 228 / direccion 227 (NOP)
"1111000000", -- linea 229 / direccion 228 (NOP)
"1111000000", -- linea 230 / direccion 229 (NOP)
"1111000000", -- linea 231 / direccion 230 (NOP)
"1111000000", -- linea 232 / direccion 231 (NOP)
"1111000000", -- linea 233 / direccion 232 (NOP)
"1111000000", -- linea 234 / direccion 233 (NOP)
"1111000000", -- linea 235 / direccion 234 (NOP)
"1111000000", -- linea 236 / direccion 235 (NOP)
"1111000000", -- linea 237 / direccion 236 (NOP)
"1111000000", -- linea 238 / direccion 237 (NOP)
"1111000000", -- linea 239 / direccion 238 (NOP)
"1111000000", -- linea 240 / direccion 239 (NOP)
"1111000000", -- linea 241 / direccion 240 (NOP)
"1111000000", -- linea 242 / direccion 241 (NOP)
"1111000000", -- linea 243 / direccion 242 (NOP)
"1111000000", -- linea 244 / direccion 243 (NOP)
"1111000000", -- linea 245 / direccion 244 (NOP)
"1111000000", -- linea 246 / direccion 245 (NOP)
"1111000000", -- linea 247 / direccion 246 (NOP)
"1111000000", -- linea 248 / direccion 247 (NOP)
"1111000000", -- linea 249 / direccion 248 (NOP)
"1111000000", -- linea 250 / direccion 249 (NOP)
"1111000000", -- linea 251 / direccion 250 (NOP)
"1111000000", -- linea 252 / direccion 251 (NOP)
"1111000000", -- linea 253 / direccion 252 (NOP)
"1111000000", -- linea 254 / direccion 253 (NOP)
"1111000000", -- linea 255 / direccion 254 (NOP)
"1111000000", -- linea 256 / direccion 255 (NOP)
"1111000000", -- linea 257 / direccion 256 (NOP)
"1111000000", -- linea 258 / direccion 257 (NOP)
"1111000000", -- linea 259 / direccion 258 (NOP)
"1111000000", -- linea 260 / direccion 259 (NOP)
"1111000000", -- linea 261 / direccion 260 (NOP)
"1111000000", -- linea 262 / direccion 261 (NOP)
"1111000000", -- linea 263 / direccion 262 (NOP)
"1111000000", -- linea 264 / direccion 263 (NOP)
"1111000000", -- linea 265 / direccion 264 (NOP)
"1111000000", -- linea 266 / direccion 265 (NOP)
"1111000000", -- linea 267 / direccion 266 (NOP)
"1111000000", -- linea 268 / direccion 267 (NOP)
"1111000000", -- linea 269 / direccion 268 (NOP)
"1111000000", -- linea 270 / direccion 269 (NOP)
"1111000000", -- linea 271 / direccion 270 (NOP)
"1111000000", -- linea 272 / direccion 271 (NOP)
"1111000000", -- linea 273 / direccion 272 (NOP)
"1111000000", -- linea 274 / direccion 273 (NOP)
"1111000000", -- linea 275 / direccion 274 (NOP)
"1111000000", -- linea 276 / direccion 275 (NOP)
"1111000000", -- linea 277 / direccion 276 (NOP)
"1111000000", -- linea 278 / direccion 277 (NOP)
"1111000000", -- linea 279 / direccion 278 (NOP)
"1111000000", -- linea 280 / direccion 279 (NOP)
"1111000000", -- linea 281 / direccion 280 (NOP)
"1111000000", -- linea 282 / direccion 281 (NOP)
"1111000000", -- linea 283 / direccion 282 (NOP)
"1111000000", -- linea 284 / direccion 283 (NOP)
"1111000000", -- linea 285 / direccion 284 (NOP)
"1111000000", -- linea 286 / direccion 285 (NOP)
"1111000000", -- linea 287 / direccion 286 (NOP)
"1111000000", -- linea 288 / direccion 287 (NOP)
"1111000000", -- linea 289 / direccion 288 (NOP)
"1111000000", -- linea 290 / direccion 289 (NOP)
"1111000000", -- linea 291 / direccion 290 (NOP)
"1111000000", -- linea 292 / direccion 291 (NOP)
"1111000000", -- linea 293 / direccion 292 (NOP)
"1111000000", -- linea 294 / direccion 293 (NOP)
"1111000000", -- linea 295 / direccion 294 (NOP)
"1111000000", -- linea 296 / direccion 295 (NOP)
"1111000000", -- linea 297 / direccion 296 (NOP)
"1111000000", -- linea 298 / direccion 297 (NOP)
"1111000000", -- linea 299 / direccion 298 (NOP)
"1111000000", -- linea 300 / direccion 299 (NOP)
"1111000000", -- linea 301 / direccion 300 (NOP)
"1111000000", -- linea 302 / direccion 301 (NOP)
"1111000000", -- linea 303 / direccion 302 (NOP)
"1111000000", -- linea 304 / direccion 303 (NOP)
"1111000000", -- linea 305 / direccion 304 (NOP)
"1111000000", -- linea 306 / direccion 305 (NOP)
"1111000000", -- linea 307 / direccion 306 (NOP)
"1111000000", -- linea 308 / direccion 307 (NOP)
"1111000000", -- linea 309 / direccion 308 (NOP)
"1111000000", -- linea 310 / direccion 309 (NOP)
"1111000000", -- linea 311 / direccion 310 (NOP)
"1111000000", -- linea 312 / direccion 311 (NOP)
"1111000000", -- linea 313 / direccion 312 (NOP)
"1111000000", -- linea 314 / direccion 313 (NOP)
"1111000000", -- linea 315 / direccion 314 (NOP)
"1111000000", -- linea 316 / direccion 315 (NOP)
"1111000000", -- linea 317 / direccion 316 (NOP)
"1111000000", -- linea 318 / direccion 317 (NOP)
"1111000000", -- linea 319 / direccion 318 (NOP)
"1111000000", -- linea 320 / direccion 319 (NOP)
"1111000000", -- linea 321 / direccion 320 (NOP)
"1111000000", -- linea 322 / direccion 321 (NOP)
"1111000000", -- linea 323 / direccion 322 (NOP)
"1111000000", -- linea 324 / direccion 323 (NOP)
"1111000000", -- linea 325 / direccion 324 (NOP)
"1111000000", -- linea 326 / direccion 325 (NOP)
"1111000000", -- linea 327 / direccion 326 (NOP)
"1111000000", -- linea 328 / direccion 327 (NOP)
"1111000000", -- linea 329 / direccion 328 (NOP)
"1111000000", -- linea 330 / direccion 329 (NOP)
"1111000000", -- linea 331 / direccion 330 (NOP)
"1111000000", -- linea 332 / direccion 331 (NOP)
"1111000000", -- linea 333 / direccion 332 (NOP)
"1111000000", -- linea 334 / direccion 333 (NOP)
"1111000000", -- linea 335 / direccion 334 (NOP)
"1111000000", -- linea 336 / direccion 335 (NOP)
"1111000000", -- linea 337 / direccion 336 (NOP)
"1111000000", -- linea 338 / direccion 337 (NOP)
"1111000000", -- linea 339 / direccion 338 (NOP)
"1111000000", -- linea 340 / direccion 339 (NOP)
"1111000000", -- linea 341 / direccion 340 (NOP)
"1111000000", -- linea 342 / direccion 341 (NOP)
"1111000000", -- linea 343 / direccion 342 (NOP)
"1111000000", -- linea 344 / direccion 343 (NOP)
"1111000000", -- linea 345 / direccion 344 (NOP)
"1111000000", -- linea 346 / direccion 345 (NOP)
"1111000000", -- linea 347 / direccion 346 (NOP)
"1111000000", -- linea 348 / direccion 347 (NOP)
"1111000000", -- linea 349 / direccion 348 (NOP)
"1111000000", -- linea 350 / direccion 349 (NOP)
"1111000000", -- linea 351 / direccion 350 (NOP)
"1111000000", -- linea 352 / direccion 351 (NOP)
"1111000000", -- linea 353 / direccion 352 (NOP)
"1111000000", -- linea 354 / direccion 353 (NOP)
"1111000000", -- linea 355 / direccion 354 (NOP)
"1111000000", -- linea 356 / direccion 355 (NOP)
"1111000000", -- linea 357 / direccion 356 (NOP)
"1111000000", -- linea 358 / direccion 357 (NOP)
"1111000000", -- linea 359 / direccion 358 (NOP)
"1111000000", -- linea 360 / direccion 359 (NOP)
"1111000000", -- linea 361 / direccion 360 (NOP)
"1111000000", -- linea 362 / direccion 361 (NOP)
"1111000000", -- linea 363 / direccion 362 (NOP)
"1111000000", -- linea 364 / direccion 363 (NOP)
"1111000000", -- linea 365 / direccion 364 (NOP)
"1111000000", -- linea 366 / direccion 365 (NOP)
"1111000000", -- linea 367 / direccion 366 (NOP)
"1111000000", -- linea 368 / direccion 367 (NOP)
"1111000000", -- linea 369 / direccion 368 (NOP)
"1111000000", -- linea 370 / direccion 369 (NOP)
"1111000000", -- linea 371 / direccion 370 (NOP)
"1111000000", -- linea 372 / direccion 371 (NOP)
"1111000000", -- linea 373 / direccion 372 (NOP)
"1111000000", -- linea 374 / direccion 373 (NOP)
"1111000000", -- linea 375 / direccion 374 (NOP)
"1111000000", -- linea 376 / direccion 375 (NOP)
"1111000000", -- linea 377 / direccion 376 (NOP)
"1111000000", -- linea 378 / direccion 377 (NOP)
"1111000000", -- linea 379 / direccion 378 (NOP)
"1111000000", -- linea 380 / direccion 379 (NOP)
"1111000000", -- linea 381 / direccion 380 (NOP)
"1111000000", -- linea 382 / direccion 381 (NOP)
"1111000000", -- linea 383 / direccion 382 (NOP)
"1111000000", -- linea 384 / direccion 383 (NOP)
"1111000000", -- linea 385 / direccion 384 (NOP)
"1111000000", -- linea 386 / direccion 385 (NOP)
"1111000000", -- linea 387 / direccion 386 (NOP)
"1111000000", -- linea 388 / direccion 387 (NOP)
"1111000000", -- linea 389 / direccion 388 (NOP)
"1111000000", -- linea 390 / direccion 389 (NOP)
"1111000000", -- linea 391 / direccion 390 (NOP)
"1111000000", -- linea 392 / direccion 391 (NOP)
"1111000000", -- linea 393 / direccion 392 (NOP)
"1111000000", -- linea 394 / direccion 393 (NOP)
"1111000000", -- linea 395 / direccion 394 (NOP)
"1111000000", -- linea 396 / direccion 395 (NOP)
"1111000000", -- linea 397 / direccion 396 (NOP)
"1111000000", -- linea 398 / direccion 397 (NOP)
"1111000000", -- linea 399 / direccion 398 (NOP)
"1111000000", -- linea 400 / direccion 399 (NOP)
"1111000000", -- linea 401 / direccion 400 (NOP)
"1111000000", -- linea 402 / direccion 401 (NOP)
"1111000000", -- linea 403 / direccion 402 (NOP)
"1111000000", -- linea 404 / direccion 403 (NOP)
"1111000000", -- linea 405 / direccion 404 (NOP)
"1111000000", -- linea 406 / direccion 405 (NOP)
"1111000000", -- linea 407 / direccion 406 (NOP)
"1111000000", -- linea 408 / direccion 407 (NOP)
"1111000000", -- linea 409 / direccion 408 (NOP)
"1111000000", -- linea 410 / direccion 409 (NOP)
"1111000000", -- linea 411 / direccion 410 (NOP)
"1111000000", -- linea 412 / direccion 411 (NOP)
"1111000000", -- linea 413 / direccion 412 (NOP)
"1111000000", -- linea 414 / direccion 413 (NOP)
"1111000000", -- linea 415 / direccion 414 (NOP)
"1111000000", -- linea 416 / direccion 415 (NOP)
"1111000000", -- linea 417 / direccion 416 (NOP)
"1111000000", -- linea 418 / direccion 417 (NOP)
"1111000000", -- linea 419 / direccion 418 (NOP)
"1111000000", -- linea 420 / direccion 419 (NOP)
"1111000000", -- linea 421 / direccion 420 (NOP)
"1111000000", -- linea 422 / direccion 421 (NOP)
"1111000000", -- linea 423 / direccion 422 (NOP)
"1111000000", -- linea 424 / direccion 423 (NOP)
"1111000000", -- linea 425 / direccion 424 (NOP)
"1111000000", -- linea 426 / direccion 425 (NOP)
"1111000000", -- linea 427 / direccion 426 (NOP)
"1111000000", -- linea 428 / direccion 427 (NOP)
"1111000000", -- linea 429 / direccion 428 (NOP)
"1111000000", -- linea 430 / direccion 429 (NOP)
"1111000000", -- linea 431 / direccion 430 (NOP)
"1111000000", -- linea 432 / direccion 431 (NOP)
"1111000000", -- linea 433 / direccion 432 (NOP)
"1111000000", -- linea 434 / direccion 433 (NOP)
"1111000000", -- linea 435 / direccion 434 (NOP)
"1111000000", -- linea 436 / direccion 435 (NOP)
"1111000000", -- linea 437 / direccion 436 (NOP)
"1111000000", -- linea 438 / direccion 437 (NOP)
"1111000000", -- linea 439 / direccion 438 (NOP)
"1111000000", -- linea 440 / direccion 439 (NOP)
"1111000000", -- linea 441 / direccion 440 (NOP)
"1111000000", -- linea 442 / direccion 441 (NOP)
"1111000000", -- linea 443 / direccion 442 (NOP)
"1111000000", -- linea 444 / direccion 443 (NOP)
"1111000000", -- linea 445 / direccion 444 (NOP)
"1111000000", -- linea 446 / direccion 445 (NOP)
"1111000000", -- linea 447 / direccion 446 (NOP)
"1111000000", -- linea 448 / direccion 447 (NOP)
"1111000000", -- linea 449 / direccion 448 (NOP)
"1111000000", -- linea 450 / direccion 449 (NOP)
"1111000000", -- linea 451 / direccion 450 (NOP)
"1111000000", -- linea 452 / direccion 451 (NOP)
"1111000000", -- linea 453 / direccion 452 (NOP)
"1111000000", -- linea 454 / direccion 453 (NOP)
"1111000000", -- linea 455 / direccion 454 (NOP)
"1111000000", -- linea 456 / direccion 455 (NOP)
"1111000000", -- linea 457 / direccion 456 (NOP)
"1111000000", -- linea 458 / direccion 457 (NOP)
"1111000000", -- linea 459 / direccion 458 (NOP)
"1111000000", -- linea 460 / direccion 459 (NOP)
"1111000000", -- linea 461 / direccion 460 (NOP)
"1111000000", -- linea 462 / direccion 461 (NOP)
"1111000000", -- linea 463 / direccion 462 (NOP)
"1111000000", -- linea 464 / direccion 463 (NOP)
"1111000000", -- linea 465 / direccion 464 (NOP)
"1111000000", -- linea 466 / direccion 465 (NOP)
"1111000000", -- linea 467 / direccion 466 (NOP)
"1111000000", -- linea 468 / direccion 467 (NOP)
"1111000000", -- linea 469 / direccion 468 (NOP)
"1111000000", -- linea 470 / direccion 469 (NOP)
"1111000000", -- linea 471 / direccion 470 (NOP)
"1111000000", -- linea 472 / direccion 471 (NOP)
"1111000000", -- linea 473 / direccion 472 (NOP)
"1111000000", -- linea 474 / direccion 473 (NOP)
"1111000000", -- linea 475 / direccion 474 (NOP)
"1111000000", -- linea 476 / direccion 475 (NOP)
"1111000000", -- linea 477 / direccion 476 (NOP)
"1111000000", -- linea 478 / direccion 477 (NOP)
"1111000000", -- linea 479 / direccion 478 (NOP)
"1111000000", -- linea 480 / direccion 479 (NOP)
"1111000000", -- linea 481 / direccion 480 (NOP)
"1111000000", -- linea 482 / direccion 481 (NOP)
"1111000000", -- linea 483 / direccion 482 (NOP)
"1111000000", -- linea 484 / direccion 483 (NOP)
"1111000000", -- linea 485 / direccion 484 (NOP)
"1111000000", -- linea 486 / direccion 485 (NOP)
"1111000000", -- linea 487 / direccion 486 (NOP)
"1111000000", -- linea 488 / direccion 487 (NOP)
"1111000000", -- linea 489 / direccion 488 (NOP)
"1111000000", -- linea 490 / direccion 489 (NOP)
"1111000000", -- linea 491 / direccion 490 (NOP)
"1111000000", -- linea 492 / direccion 491 (NOP)
"1111000000", -- linea 493 / direccion 492 (NOP)
"1111000000", -- linea 494 / direccion 493 (NOP)
"1111000000", -- linea 495 / direccion 494 (NOP)
"1111000000", -- linea 496 / direccion 495 (NOP)
"1111000000", -- linea 497 / direccion 496 (NOP)
"1111000000", -- linea 498 / direccion 497 (NOP)
"1111000000", -- linea 499 / direccion 498 (NOP)
"1111000000", -- linea 500 / direccion 499 (NOP)
"1111000000", -- linea 501 / direccion 500 (NOP)
"1111000000", -- linea 502 / direccion 501 (NOP)
"1111000000", -- linea 503 / direccion 502 (NOP)
"1111000000", -- linea 504 / direccion 503 (NOP)
"1111000000", -- linea 505 / direccion 504 (NOP)
"1111000000", -- linea 506 / direccion 505 (NOP)
"1111000000", -- linea 507 / direccion 506 (NOP)
"1111000000", -- linea 508 / direccion 507 (NOP)
"1111000000", -- linea 509 / direccion 508 (NOP)
"1111000000", -- linea 510 / direccion 509 (NOP)
"1111000000", -- linea 511 / direccion 510 (NOP)
"1111000000", -- linea 512 / direccion 511 (NOP)
"1111000000", -- linea 513 / direccion 512 (NOP)
"1111000000", -- linea 514 / direccion 513 (NOP)
"1111000000", -- linea 515 / direccion 514 (NOP)
"1111000000", -- linea 516 / direccion 515 (NOP)
"1111000000", -- linea 517 / direccion 516 (NOP)
"1111000000", -- linea 518 / direccion 517 (NOP)
"1111000000", -- linea 519 / direccion 518 (NOP)
"1111000000", -- linea 520 / direccion 519 (NOP)
"1111000000", -- linea 521 / direccion 520 (NOP)
"1111000000", -- linea 522 / direccion 521 (NOP)
"1111000000", -- linea 523 / direccion 522 (NOP)
"1111000000", -- linea 524 / direccion 523 (NOP)
"1111000000", -- linea 525 / direccion 524 (NOP)
"1111000000", -- linea 526 / direccion 525 (NOP)
"1111000000", -- linea 527 / direccion 526 (NOP)
"1111000000", -- linea 528 / direccion 527 (NOP)
"1111000000", -- linea 529 / direccion 528 (NOP)
"1111000000", -- linea 530 / direccion 529 (NOP)
"1111000000", -- linea 531 / direccion 530 (NOP)
"1111000000", -- linea 532 / direccion 531 (NOP)
"1111000000", -- linea 533 / direccion 532 (NOP)
"1111000000", -- linea 534 / direccion 533 (NOP)
"1111000000", -- linea 535 / direccion 534 (NOP)
"1111000000", -- linea 536 / direccion 535 (NOP)
"1111000000", -- linea 537 / direccion 536 (NOP)
"1111000000", -- linea 538 / direccion 537 (NOP)
"1111000000", -- linea 539 / direccion 538 (NOP)
"1111000000", -- linea 540 / direccion 539 (NOP)
"1111000000", -- linea 541 / direccion 540 (NOP)
"1111000000", -- linea 542 / direccion 541 (NOP)
"1111000000", -- linea 543 / direccion 542 (NOP)
"1111000000", -- linea 544 / direccion 543 (NOP)
"1111000000", -- linea 545 / direccion 544 (NOP)
"1111000000", -- linea 546 / direccion 545 (NOP)
"1111000000", -- linea 547 / direccion 546 (NOP)
"1111000000", -- linea 548 / direccion 547 (NOP)
"1111000000", -- linea 549 / direccion 548 (NOP)
"1111000000", -- linea 550 / direccion 549 (NOP)
"1111000000", -- linea 551 / direccion 550 (NOP)
"1111000000", -- linea 552 / direccion 551 (NOP)
"1111000000", -- linea 553 / direccion 552 (NOP)
"1111000000", -- linea 554 / direccion 553 (NOP)
"1111000000", -- linea 555 / direccion 554 (NOP)
"1111000000", -- linea 556 / direccion 555 (NOP)
"1111000000", -- linea 557 / direccion 556 (NOP)
"1111000000", -- linea 558 / direccion 557 (NOP)
"1111000000", -- linea 559 / direccion 558 (NOP)
"1111000000", -- linea 560 / direccion 559 (NOP)
"1111000000", -- linea 561 / direccion 560 (NOP)
"1111000000", -- linea 562 / direccion 561 (NOP)
"1111000000", -- linea 563 / direccion 562 (NOP)
"1111000000", -- linea 564 / direccion 563 (NOP)
"1111000000", -- linea 565 / direccion 564 (NOP)
"1111000000", -- linea 566 / direccion 565 (NOP)
"1111000000", -- linea 567 / direccion 566 (NOP)
"1111000000", -- linea 568 / direccion 567 (NOP)
"1111000000", -- linea 569 / direccion 568 (NOP)
"1111000000", -- linea 570 / direccion 569 (NOP)
"1111000000", -- linea 571 / direccion 570 (NOP)
"1111000000", -- linea 572 / direccion 571 (NOP)
"1111000000", -- linea 573 / direccion 572 (NOP)
"1111000000", -- linea 574 / direccion 573 (NOP)
"1111000000", -- linea 575 / direccion 574 (NOP)
"1111000000", -- linea 576 / direccion 575 (NOP)
"1111000000", -- linea 577 / direccion 576 (NOP)
"1111000000", -- linea 578 / direccion 577 (NOP)
"1111000000", -- linea 579 / direccion 578 (NOP)
"1111000000", -- linea 580 / direccion 579 (NOP)
"1111000000", -- linea 581 / direccion 580 (NOP)
"1111000000", -- linea 582 / direccion 581 (NOP)
"1111000000", -- linea 583 / direccion 582 (NOP)
"1111000000", -- linea 584 / direccion 583 (NOP)
"1111000000", -- linea 585 / direccion 584 (NOP)
"1111000000", -- linea 586 / direccion 585 (NOP)
"1111000000", -- linea 587 / direccion 586 (NOP)
"1111000000", -- linea 588 / direccion 587 (NOP)
"1111000000", -- linea 589 / direccion 588 (NOP)
"1111000000", -- linea 590 / direccion 589 (NOP)
"1111000000", -- linea 591 / direccion 590 (NOP)
"1111000000", -- linea 592 / direccion 591 (NOP)
"1111000000", -- linea 593 / direccion 592 (NOP)
"1111000000", -- linea 594 / direccion 593 (NOP)
"1111000000", -- linea 595 / direccion 594 (NOP)
"1111000000", -- linea 596 / direccion 595 (NOP)
"1111000000", -- linea 597 / direccion 596 (NOP)
"1111000000", -- linea 598 / direccion 597 (NOP)
"1111000000", -- linea 599 / direccion 598 (NOP)
"1111000000", -- linea 600 / direccion 599 (NOP)
"1111000000", -- linea 601 / direccion 600 (NOP)
"1111000000", -- linea 602 / direccion 601 (NOP)
"1111000000", -- linea 603 / direccion 602 (NOP)
"1111000000", -- linea 604 / direccion 603 (NOP)
"1111000000", -- linea 605 / direccion 604 (NOP)
"1111000000", -- linea 606 / direccion 605 (NOP)
"1111000000", -- linea 607 / direccion 606 (NOP)
"1111000000", -- linea 608 / direccion 607 (NOP)
"1111000000", -- linea 609 / direccion 608 (NOP)
"1111000000", -- linea 610 / direccion 609 (NOP)
"1111000000", -- linea 611 / direccion 610 (NOP)
"1111000000", -- linea 612 / direccion 611 (NOP)
"1111000000", -- linea 613 / direccion 612 (NOP)
"1111000000", -- linea 614 / direccion 613 (NOP)
"1111000000", -- linea 615 / direccion 614 (NOP)
"1111000000", -- linea 616 / direccion 615 (NOP)
"1111000000", -- linea 617 / direccion 616 (NOP)
"1111000000", -- linea 618 / direccion 617 (NOP)
"1111000000", -- linea 619 / direccion 618 (NOP)
"1111000000", -- linea 620 / direccion 619 (NOP)
"1111000000", -- linea 621 / direccion 620 (NOP)
"1111000000", -- linea 622 / direccion 621 (NOP)
"1111000000", -- linea 623 / direccion 622 (NOP)
"1111000000", -- linea 624 / direccion 623 (NOP)
"1111000000", -- linea 625 / direccion 624 (NOP)
"1111000000", -- linea 626 / direccion 625 (NOP)
"1111000000", -- linea 627 / direccion 626 (NOP)
"1111000000", -- linea 628 / direccion 627 (NOP)
"1111000000", -- linea 629 / direccion 628 (NOP)
"1111000000", -- linea 630 / direccion 629 (NOP)
"1111000000", -- linea 631 / direccion 630 (NOP)
"1111000000", -- linea 632 / direccion 631 (NOP)
"1111000000", -- linea 633 / direccion 632 (NOP)
"1111000000", -- linea 634 / direccion 633 (NOP)
"1111000000", -- linea 635 / direccion 634 (NOP)
"1111000000", -- linea 636 / direccion 635 (NOP)
"1111000000", -- linea 637 / direccion 636 (NOP)
"1111000000", -- linea 638 / direccion 637 (NOP)
"1111000000", -- linea 639 / direccion 638 (NOP)
"1111000000", -- linea 640 / direccion 639 (NOP)
"1111000000", -- linea 641 / direccion 640 (NOP)
"1111000000", -- linea 642 / direccion 641 (NOP)
"1111000000", -- linea 643 / direccion 642 (NOP)
"1111000000", -- linea 644 / direccion 643 (NOP)
"1111000000", -- linea 645 / direccion 644 (NOP)
"1111000000", -- linea 646 / direccion 645 (NOP)
"1111000000", -- linea 647 / direccion 646 (NOP)
"1111000000", -- linea 648 / direccion 647 (NOP)
"1111000000", -- linea 649 / direccion 648 (NOP)
"1111000000", -- linea 650 / direccion 649 (NOP)
"1111000000", -- linea 651 / direccion 650 (NOP)
"1111000000", -- linea 652 / direccion 651 (NOP)
"1111000000", -- linea 653 / direccion 652 (NOP)
"1111000000", -- linea 654 / direccion 653 (NOP)
"1111000000", -- linea 655 / direccion 654 (NOP)
"1111000000", -- linea 656 / direccion 655 (NOP)
"1111000000", -- linea 657 / direccion 656 (NOP)
"1111000000", -- linea 658 / direccion 657 (NOP)
"1111000000", -- linea 659 / direccion 658 (NOP)
"1111000000", -- linea 660 / direccion 659 (NOP)
"1111000000", -- linea 661 / direccion 660 (NOP)
"1111000000", -- linea 662 / direccion 661 (NOP)
"1111000000", -- linea 663 / direccion 662 (NOP)
"1111000000", -- linea 664 / direccion 663 (NOP)
"1111000000", -- linea 665 / direccion 664 (NOP)
"1111000000", -- linea 666 / direccion 665 (NOP)
"1111000000", -- linea 667 / direccion 666 (NOP)
"1111000000", -- linea 668 / direccion 667 (NOP)
"1111000000", -- linea 669 / direccion 668 (NOP)
"1111000000", -- linea 670 / direccion 669 (NOP)
"1111000000", -- linea 671 / direccion 670 (NOP)
"1111000000", -- linea 672 / direccion 671 (NOP)
"1111000000", -- linea 673 / direccion 672 (NOP)
"1111000000", -- linea 674 / direccion 673 (NOP)
"1111000000", -- linea 675 / direccion 674 (NOP)
"1111000000", -- linea 676 / direccion 675 (NOP)
"1111000000", -- linea 677 / direccion 676 (NOP)
"1111000000", -- linea 678 / direccion 677 (NOP)
"1111000000", -- linea 679 / direccion 678 (NOP)
"1111000000", -- linea 680 / direccion 679 (NOP)
"1111000000", -- linea 681 / direccion 680 (NOP)
"1111000000", -- linea 682 / direccion 681 (NOP)
"1111000000", -- linea 683 / direccion 682 (NOP)
"1111000000", -- linea 684 / direccion 683 (NOP)
"1111000000", -- linea 685 / direccion 684 (NOP)
"1111000000", -- linea 686 / direccion 685 (NOP)
"1111000000", -- linea 687 / direccion 686 (NOP)
"1111000000", -- linea 688 / direccion 687 (NOP)
"1111000000", -- linea 689 / direccion 688 (NOP)
"1111000000", -- linea 690 / direccion 689 (NOP)
"1111000000", -- linea 691 / direccion 690 (NOP)
"1111000000", -- linea 692 / direccion 691 (NOP)
"1111000000", -- linea 693 / direccion 692 (NOP)
"1111000000", -- linea 694 / direccion 693 (NOP)
"1111000000", -- linea 695 / direccion 694 (NOP)
"1111000000", -- linea 696 / direccion 695 (NOP)
"1111000000", -- linea 697 / direccion 696 (NOP)
"1111000000", -- linea 698 / direccion 697 (NOP)
"1111000000", -- linea 699 / direccion 698 (NOP)
"1111000000", -- linea 700 / direccion 699 (NOP)
"1111000000", -- linea 701 / direccion 700 (NOP)
"1111000000", -- linea 702 / direccion 701 (NOP)
"1111000000", -- linea 703 / direccion 702 (NOP)
"1111000000", -- linea 704 / direccion 703 (NOP)
"1111000000", -- linea 705 / direccion 704 (NOP)
"1111000000", -- linea 706 / direccion 705 (NOP)
"1111000000", -- linea 707 / direccion 706 (NOP)
"1111000000", -- linea 708 / direccion 707 (NOP)
"1111000000", -- linea 709 / direccion 708 (NOP)
"1111000000", -- linea 710 / direccion 709 (NOP)
"1111000000", -- linea 711 / direccion 710 (NOP)
"1111000000", -- linea 712 / direccion 711 (NOP)
"1111000000", -- linea 713 / direccion 712 (NOP)
"1111000000", -- linea 714 / direccion 713 (NOP)
"1111000000", -- linea 715 / direccion 714 (NOP)
"1111000000", -- linea 716 / direccion 715 (NOP)
"1111000000", -- linea 717 / direccion 716 (NOP)
"1111000000", -- linea 718 / direccion 717 (NOP)
"1111000000", -- linea 719 / direccion 718 (NOP)
"1111000000", -- linea 720 / direccion 719 (NOP)
"1111000000", -- linea 721 / direccion 720 (NOP)
"1111000000", -- linea 722 / direccion 721 (NOP)
"1111000000", -- linea 723 / direccion 722 (NOP)
"1111000000", -- linea 724 / direccion 723 (NOP)
"1111000000", -- linea 725 / direccion 724 (NOP)
"1111000000", -- linea 726 / direccion 725 (NOP)
"1111000000", -- linea 727 / direccion 726 (NOP)
"1111000000", -- linea 728 / direccion 727 (NOP)
"1111000000", -- linea 729 / direccion 728 (NOP)
"1111000000", -- linea 730 / direccion 729 (NOP)
"1111000000", -- linea 731 / direccion 730 (NOP)
"1111000000", -- linea 732 / direccion 731 (NOP)
"1111000000", -- linea 733 / direccion 732 (NOP)
"1111000000", -- linea 734 / direccion 733 (NOP)
"1111000000", -- linea 735 / direccion 734 (NOP)
"1111000000", -- linea 736 / direccion 735 (NOP)
"1111000000", -- linea 737 / direccion 736 (NOP)
"1111000000", -- linea 738 / direccion 737 (NOP)
"1111000000", -- linea 739 / direccion 738 (NOP)
"1111000000", -- linea 740 / direccion 739 (NOP)
"1111000000", -- linea 741 / direccion 740 (NOP)
"1111000000", -- linea 742 / direccion 741 (NOP)
"1111000000", -- linea 743 / direccion 742 (NOP)
"1111000000", -- linea 744 / direccion 743 (NOP)
"1111000000", -- linea 745 / direccion 744 (NOP)
"1111000000", -- linea 746 / direccion 745 (NOP)
"1111000000", -- linea 747 / direccion 746 (NOP)
"1111000000", -- linea 748 / direccion 747 (NOP)
"1111000000", -- linea 749 / direccion 748 (NOP)
"1111000000", -- linea 750 / direccion 749 (NOP)
"1111000000", -- linea 751 / direccion 750 (NOP)
"1111000000", -- linea 752 / direccion 751 (NOP)
"1111000000", -- linea 753 / direccion 752 (NOP)
"1111000000", -- linea 754 / direccion 753 (NOP)
"1111000000", -- linea 755 / direccion 754 (NOP)
"1111000000", -- linea 756 / direccion 755 (NOP)
"1111000000", -- linea 757 / direccion 756 (NOP)
"1111000000", -- linea 758 / direccion 757 (NOP)
"1111000000", -- linea 759 / direccion 758 (NOP)
"1111000000", -- linea 760 / direccion 759 (NOP)
"1111000000", -- linea 761 / direccion 760 (NOP)
"1111000000", -- linea 762 / direccion 761 (NOP)
"1111000000", -- linea 763 / direccion 762 (NOP)
"1111000000", -- linea 764 / direccion 763 (NOP)
"1111000000", -- linea 765 / direccion 764 (NOP)
"1111000000", -- linea 766 / direccion 765 (NOP)
"1111000000", -- linea 767 / direccion 766 (NOP)
"1111000000", -- linea 768 / direccion 767 (NOP)
"1111000000", -- linea 769 / direccion 768 (NOP)
"1111000000", -- linea 770 / direccion 769 (NOP)
"1111000000", -- linea 771 / direccion 770 (NOP)
"1111000000", -- linea 772 / direccion 771 (NOP)
"1111000000", -- linea 773 / direccion 772 (NOP)
"1111000000", -- linea 774 / direccion 773 (NOP)
"1111000000", -- linea 775 / direccion 774 (NOP)
"1111000000", -- linea 776 / direccion 775 (NOP)
"1111000000", -- linea 777 / direccion 776 (NOP)
"1111000000", -- linea 778 / direccion 777 (NOP)
"1111000000", -- linea 779 / direccion 778 (NOP)
"1111000000", -- linea 780 / direccion 779 (NOP)
"1111000000", -- linea 781 / direccion 780 (NOP)
"1111000000", -- linea 782 / direccion 781 (NOP)
"1111000000", -- linea 783 / direccion 782 (NOP)
"1111000000", -- linea 784 / direccion 783 (NOP)
"1111000000", -- linea 785 / direccion 784 (NOP)
"1111000000", -- linea 786 / direccion 785 (NOP)
"1111000000", -- linea 787 / direccion 786 (NOP)
"1111000000", -- linea 788 / direccion 787 (NOP)
"1111000000", -- linea 789 / direccion 788 (NOP)
"1111000000", -- linea 790 / direccion 789 (NOP)
"1111000000", -- linea 791 / direccion 790 (NOP)
"1111000000", -- linea 792 / direccion 791 (NOP)
"1111000000", -- linea 793 / direccion 792 (NOP)
"1111000000", -- linea 794 / direccion 793 (NOP)
"1111000000", -- linea 795 / direccion 794 (NOP)
"1111000000", -- linea 796 / direccion 795 (NOP)
"1111000000", -- linea 797 / direccion 796 (NOP)
"1111000000", -- linea 798 / direccion 797 (NOP)
"1111000000", -- linea 799 / direccion 798 (NOP)
"1111000000", -- linea 800 / direccion 799 (NOP)
"1111000000", -- linea 801 / direccion 800 (NOP)
"1111000000", -- linea 802 / direccion 801 (NOP)
"1111000000", -- linea 803 / direccion 802 (NOP)
"1111000000", -- linea 804 / direccion 803 (NOP)
"1111000000", -- linea 805 / direccion 804 (NOP)
"1111000000", -- linea 806 / direccion 805 (NOP)
"1111000000", -- linea 807 / direccion 806 (NOP)
"1111000000", -- linea 808 / direccion 807 (NOP)
"1111000000", -- linea 809 / direccion 808 (NOP)
"1111000000", -- linea 810 / direccion 809 (NOP)
"1111000000", -- linea 811 / direccion 810 (NOP)
"1111000000", -- linea 812 / direccion 811 (NOP)
"1111000000", -- linea 813 / direccion 812 (NOP)
"1111000000", -- linea 814 / direccion 813 (NOP)
"1111000000", -- linea 815 / direccion 814 (NOP)
"1111000000", -- linea 816 / direccion 815 (NOP)
"1111000000", -- linea 817 / direccion 816 (NOP)
"1111000000", -- linea 818 / direccion 817 (NOP)
"1111000000", -- linea 819 / direccion 818 (NOP)
"1111000000", -- linea 820 / direccion 819 (NOP)
"1111000000", -- linea 821 / direccion 820 (NOP)
"1111000000", -- linea 822 / direccion 821 (NOP)
"1111000000", -- linea 823 / direccion 822 (NOP)
"1111000000", -- linea 824 / direccion 823 (NOP)
"1111000000", -- linea 825 / direccion 824 (NOP)
"1111000000", -- linea 826 / direccion 825 (NOP)
"1111000000", -- linea 827 / direccion 826 (NOP)
"1111000000", -- linea 828 / direccion 827 (NOP)
"1111000000", -- linea 829 / direccion 828 (NOP)
"1111000000", -- linea 830 / direccion 829 (NOP)
"1111000000", -- linea 831 / direccion 830 (NOP)
"1111000000", -- linea 832 / direccion 831 (NOP)
"1111000000", -- linea 833 / direccion 832 (NOP)
"1111000000", -- linea 834 / direccion 833 (NOP)
"1111000000", -- linea 835 / direccion 834 (NOP)
"1111000000", -- linea 836 / direccion 835 (NOP)
"1111000000", -- linea 837 / direccion 836 (NOP)
"1111000000", -- linea 838 / direccion 837 (NOP)
"1111000000", -- linea 839 / direccion 838 (NOP)
"1111000000", -- linea 840 / direccion 839 (NOP)
"1111000000", -- linea 841 / direccion 840 (NOP)
"1111000000", -- linea 842 / direccion 841 (NOP)
"1111000000", -- linea 843 / direccion 842 (NOP)
"1111000000", -- linea 844 / direccion 843 (NOP)
"1111000000", -- linea 845 / direccion 844 (NOP)
"1111000000", -- linea 846 / direccion 845 (NOP)
"1111000000", -- linea 847 / direccion 846 (NOP)
"1111000000", -- linea 848 / direccion 847 (NOP)
"1111000000", -- linea 849 / direccion 848 (NOP)
"1111000000", -- linea 850 / direccion 849 (NOP)
"1111000000", -- linea 851 / direccion 850 (NOP)
"1111000000", -- linea 852 / direccion 851 (NOP)
"1111000000", -- linea 853 / direccion 852 (NOP)
"1111000000", -- linea 854 / direccion 853 (NOP)
"1111000000", -- linea 855 / direccion 854 (NOP)
"1111000000", -- linea 856 / direccion 855 (NOP)
"1111000000", -- linea 857 / direccion 856 (NOP)
"1111000000", -- linea 858 / direccion 857 (NOP)
"1111000000", -- linea 859 / direccion 858 (NOP)
"1111000000", -- linea 860 / direccion 859 (NOP)
"1111000000", -- linea 861 / direccion 860 (NOP)
"1111000000", -- linea 862 / direccion 861 (NOP)
"1111000000", -- linea 863 / direccion 862 (NOP)
"1111000000", -- linea 864 / direccion 863 (NOP)
"1111000000", -- linea 865 / direccion 864 (NOP)
"1111000000", -- linea 866 / direccion 865 (NOP)
"1111000000", -- linea 867 / direccion 866 (NOP)
"1111000000", -- linea 868 / direccion 867 (NOP)
"1111000000", -- linea 869 / direccion 868 (NOP)
"1111000000", -- linea 870 / direccion 869 (NOP)
"1111000000", -- linea 871 / direccion 870 (NOP)
"1111000000", -- linea 872 / direccion 871 (NOP)
"1111000000", -- linea 873 / direccion 872 (NOP)
"1111000000", -- linea 874 / direccion 873 (NOP)
"1111000000", -- linea 875 / direccion 874 (NOP)
"1111000000", -- linea 876 / direccion 875 (NOP)
"1111000000", -- linea 877 / direccion 876 (NOP)
"1111000000", -- linea 878 / direccion 877 (NOP)
"1111000000", -- linea 879 / direccion 878 (NOP)
"1111000000", -- linea 880 / direccion 879 (NOP)
"1111000000", -- linea 881 / direccion 880 (NOP)
"1111000000", -- linea 882 / direccion 881 (NOP)
"1111000000", -- linea 883 / direccion 882 (NOP)
"1111000000", -- linea 884 / direccion 883 (NOP)
"1111000000", -- linea 885 / direccion 884 (NOP)
"1111000000", -- linea 886 / direccion 885 (NOP)
"1111000000", -- linea 887 / direccion 886 (NOP)
"1111000000", -- linea 888 / direccion 887 (NOP)
"1111000000", -- linea 889 / direccion 888 (NOP)
"1111000000", -- linea 890 / direccion 889 (NOP)
"1111000000", -- linea 891 / direccion 890 (NOP)
"1111000000", -- linea 892 / direccion 891 (NOP)
"1111000000", -- linea 893 / direccion 892 (NOP)
"1111000000", -- linea 894 / direccion 893 (NOP)
"1111000000", -- linea 895 / direccion 894 (NOP)
"1111000000", -- linea 896 / direccion 895 (NOP)
"1111000000", -- linea 897 / direccion 896 (NOP)
"1111000000", -- linea 898 / direccion 897 (NOP)
"1111000000", -- linea 899 / direccion 898 (NOP)
"1111000000", -- linea 900 / direccion 899 (NOP)
"1111000000", -- linea 901 / direccion 900 (NOP)
"1111000000", -- linea 902 / direccion 901 (NOP)
"1111000000", -- linea 903 / direccion 902 (NOP)
"1111000000", -- linea 904 / direccion 903 (NOP)
"1111000000", -- linea 905 / direccion 904 (NOP)
"1111000000", -- linea 906 / direccion 905 (NOP)
"1111000000", -- linea 907 / direccion 906 (NOP)
"1111000000", -- linea 908 / direccion 907 (NOP)
"1111000000", -- linea 909 / direccion 908 (NOP)
"1111000000", -- linea 910 / direccion 909 (NOP)
"1111000000", -- linea 911 / direccion 910 (NOP)
"1111000000", -- linea 912 / direccion 911 (NOP)
"1111000000", -- linea 913 / direccion 912 (NOP)
"1111000000", -- linea 914 / direccion 913 (NOP)
"1111000000", -- linea 915 / direccion 914 (NOP)
"1111000000", -- linea 916 / direccion 915 (NOP)
"1111000000", -- linea 917 / direccion 916 (NOP)
"1111000000", -- linea 918 / direccion 917 (NOP)
"1111000000", -- linea 919 / direccion 918 (NOP)
"1111000000", -- linea 920 / direccion 919 (NOP)
"1111000000", -- linea 921 / direccion 920 (NOP)
"1111000000", -- linea 922 / direccion 921 (NOP)
"1111000000", -- linea 923 / direccion 922 (NOP)
"1111000000", -- linea 924 / direccion 923 (NOP)
"1111000000", -- linea 925 / direccion 924 (NOP)
"1111000000", -- linea 926 / direccion 925 (NOP)
"1111000000", -- linea 927 / direccion 926 (NOP)
"1111000000", -- linea 928 / direccion 927 (NOP)
"1111000000", -- linea 929 / direccion 928 (NOP)
"1111000000", -- linea 930 / direccion 929 (NOP)
"1111000000", -- linea 931 / direccion 930 (NOP)
"1111000000", -- linea 932 / direccion 931 (NOP)
"1111000000", -- linea 933 / direccion 932 (NOP)
"1111000000", -- linea 934 / direccion 933 (NOP)
"1111000000", -- linea 935 / direccion 934 (NOP)
"1111000000", -- linea 936 / direccion 935 (NOP)
"1111000000", -- linea 937 / direccion 936 (NOP)
"1111000000", -- linea 938 / direccion 937 (NOP)
"1111000000", -- linea 939 / direccion 938 (NOP)
"1111000000", -- linea 940 / direccion 939 (NOP)
"1111000000", -- linea 941 / direccion 940 (NOP)
"1111000000", -- linea 942 / direccion 941 (NOP)
"1111000000", -- linea 943 / direccion 942 (NOP)
"1111000000", -- linea 944 / direccion 943 (NOP)
"1111000000", -- linea 945 / direccion 944 (NOP)
"1111000000", -- linea 946 / direccion 945 (NOP)
"1111000000", -- linea 947 / direccion 946 (NOP)
"1111000000", -- linea 948 / direccion 947 (NOP)
"1111000000", -- linea 949 / direccion 948 (NOP)
"1111000000", -- linea 950 / direccion 949 (NOP)
"1111000000", -- linea 951 / direccion 950 (NOP)
"1111000000", -- linea 952 / direccion 951 (NOP)
"1111000000", -- linea 953 / direccion 952 (NOP)
"1111000000", -- linea 954 / direccion 953 (NOP)
"1111000000", -- linea 955 / direccion 954 (NOP)
"1111000000", -- linea 956 / direccion 955 (NOP)
"1111000000", -- linea 957 / direccion 956 (NOP)
"1111000000", -- linea 958 / direccion 957 (NOP)
"1111000000", -- linea 959 / direccion 958 (NOP)
"1111000000", -- linea 960 / direccion 959 (NOP)
"1111000000", -- linea 961 / direccion 960 (NOP)
"1111000000", -- linea 962 / direccion 961 (NOP)
"1111000000", -- linea 963 / direccion 962 (NOP)
"1111000000", -- linea 964 / direccion 963 (NOP)
"1111000000", -- linea 965 / direccion 964 (NOP)
"1111000000", -- linea 966 / direccion 965 (NOP)
"1111000000", -- linea 967 / direccion 966 (NOP)
"1111000000", -- linea 968 / direccion 967 (NOP)
"1111000000", -- linea 969 / direccion 968 (NOP)
"1111000000", -- linea 970 / direccion 969 (NOP)
"1111000000", -- linea 971 / direccion 970 (NOP)
"1111000000", -- linea 972 / direccion 971 (NOP)
"1111000000", -- linea 973 / direccion 972 (NOP)
"1111000000", -- linea 974 / direccion 973 (NOP)
"1111000000", -- linea 975 / direccion 974 (NOP)
"1111000000", -- linea 976 / direccion 975 (NOP)
"1111000000", -- linea 977 / direccion 976 (NOP)
"1111000000", -- linea 978 / direccion 977 (NOP)
"1111000000", -- linea 979 / direccion 978 (NOP)
"1111000000", -- linea 980 / direccion 979 (NOP)
"1111000000", -- linea 981 / direccion 980 (NOP)
"1111000000", -- linea 982 / direccion 981 (NOP)
"1111000000", -- linea 983 / direccion 982 (NOP)
"1111000000", -- linea 984 / direccion 983 (NOP)
"1111000000", -- linea 985 / direccion 984 (NOP)
"1111000000", -- linea 986 / direccion 985 (NOP)
"1111000000", -- linea 987 / direccion 986 (NOP)
"1111000000", -- linea 988 / direccion 987 (NOP)
"1111000000", -- linea 989 / direccion 988 (NOP)
"1111000000", -- linea 990 / direccion 989 (NOP)
"1111000000", -- linea 991 / direccion 990 (NOP)
"1111000000", -- linea 992 / direccion 991 (NOP)
"1111000000", -- linea 993 / direccion 992 (NOP)
"1111000000", -- linea 994 / direccion 993 (NOP)
"1111000000", -- linea 995 / direccion 994 (NOP)
"1111000000", -- linea 996 / direccion 995 (NOP)
"1111000000", -- linea 997 / direccion 996 (NOP)
"1111000000", -- linea 998 / direccion 997 (NOP)
"1111000000", -- linea 999 / direccion 998 (NOP)
"1111000000", -- linea 1000 / direccion 999 (NOP)
"1111000000", -- linea 1001 / direccion 1000 (NOP)
"1111000000", -- linea 1002 / direccion 1001 (NOP)
"1111000000", -- linea 1003 / direccion 1002 (NOP)
"1111000000", -- linea 1004 / direccion 1003 (NOP)
"1111000000", -- linea 1005 / direccion 1004 (NOP)
"1111000000", -- linea 1006 / direccion 1005 (NOP)
"1111000000", -- linea 1007 / direccion 1006 (NOP)
"1111000000", -- linea 1008 / direccion 1007 (NOP)
"1111000000", -- linea 1009 / direccion 1008 (NOP)
"1111000000", -- linea 1010 / direccion 1009 (NOP)
"1111000000", -- linea 1011 / direccion 1010 (NOP)
"1111000000", -- linea 1012 / direccion 1011 (NOP)
"1111000000", -- linea 1013 / direccion 1012 (NOP)
"1111000000", -- linea 1014 / direccion 1013 (NOP)
"1111000000", -- linea 1015 / direccion 1014 (NOP)
"1111000000", -- linea 1016 / direccion 1015 (NOP)
"1111000000", -- linea 1017 / direccion 1016 (NOP)
"1111000000", -- linea 1018 / direccion 1017 (NOP)
"1111000000", -- linea 1019 / direccion 1018 (NOP)
"1111000000", -- linea 1020 / direccion 1019 (NOP)
"1111000000", -- linea 1021 / direccion 1020 (NOP)
"1111000000", -- linea 1022 / direccion 1021 (NOP)
"1111000000", -- linea 1023 / direccion 1022 (NOP)
"1111000000", -- linea 1024 / direccion 1023 (NOP)
		others => (others => '0')
	);

begin

	data <= ROM(to_integer(unsigned(addr)));

end arq1;
